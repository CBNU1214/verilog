/*
  Author: Jung Gyu Min.
  Affiliation: EPIC Lab, POSTECH EE.
  Description: read-only memory containing hex-code of bios program.
*/

module bios_mem_print (
    input clk,
    input ena,
    input rst,
    input [10:0] addra,
    output reg [31:0] douta,
    input enb,
    input [10:0] addrb,
    output reg [31:0] doutb
);
    wire [31:0] mem [2048-1:0];
    always @(posedge clk) begin
        if (rst) begin
            douta <= 32'b0;
        end
        else if (ena) begin
            douta <= mem[addra];
        end
    end

    always @(posedge clk) begin
        if (rst) begin
            doutb <= 32'b0;
        end
        else if (enb) begin
            doutb <= mem[addrb];
        end
    end
    
assign	mem[11'd0]	=	32'h	10010137	;
assign	mem[11'd1]	=	32'h	ff010113	;
assign	mem[11'd2]	=	32'h	1f0000ef	;
assign	mem[11'd3]	=	32'h	fd010113	;
assign	mem[11'd4]	=	32'h	02112623	;
assign	mem[11'd5]	=	32'h	02812423	;
assign	mem[11'd6]	=	32'h	02912223	;
assign	mem[11'd7]	=	32'h	03010413	;
assign	mem[11'd8]	=	32'h	fca42e23	;
assign	mem[11'd9]	=	32'h	fcb42c23	;
assign	mem[11'd10]	=	32'h	fe042623	;
assign	mem[11'd11]	=	32'h	0280006f	;
assign	mem[11'd12]	=	32'h	fdc42703	;
assign	mem[11'd13]	=	32'h	fec42783	;
assign	mem[11'd14]	=	32'h	00f704b3	;
assign	mem[11'd15]	=	32'h	7f9000ef	;
assign	mem[11'd16]	=	32'h	00050793	;
assign	mem[11'd17]	=	32'h	00f48023	;
assign	mem[11'd18]	=	32'h	fec42783	;
assign	mem[11'd19]	=	32'h	00178793	;
assign	mem[11'd20]	=	32'h	fef42623	;
assign	mem[11'd21]	=	32'h	fec42703	;
assign	mem[11'd22]	=	32'h	fd842783	;
assign	mem[11'd23]	=	32'h	fcf76ae3	;
assign	mem[11'd24]	=	32'h	fdc42703	;
assign	mem[11'd25]	=	32'h	fd842783	;
assign	mem[11'd26]	=	32'h	00f707b3	;
assign	mem[11'd27]	=	32'h	00078023	;
assign	mem[11'd28]	=	32'h	fdc42783	;
assign	mem[11'd29]	=	32'h	00078513	;
assign	mem[11'd30]	=	32'h	02c12083	;
assign	mem[11'd31]	=	32'h	02812403	;
assign	mem[11'd32]	=	32'h	02412483	;
assign	mem[11'd33]	=	32'h	03010113	;
assign	mem[11'd34]	=	32'h	00008067	;
assign	mem[11'd35]	=	32'h	fd010113	;
assign	mem[11'd36]	=	32'h	02112623	;
assign	mem[11'd37]	=	32'h	02812423	;
assign	mem[11'd38]	=	32'h	03010413	;
assign	mem[11'd39]	=	32'h	fca42e23	;
assign	mem[11'd40]	=	32'h	fcb42c23	;
assign	mem[11'd41]	=	32'h	fcc42a23	;
assign	mem[11'd42]	=	32'h	fe042623	;
assign	mem[11'd43]	=	32'h	0880006f	;
assign	mem[11'd44]	=	32'h	785000ef	;
assign	mem[11'd45]	=	32'h	00050793	;
assign	mem[11'd46]	=	32'h	fef403a3	;
assign	mem[11'd47]	=	32'h	fe042423	;
assign	mem[11'd48]	=	32'h	0400006f	;
assign	mem[11'd49]	=	32'h	fd442703	;
assign	mem[11'd50]	=	32'h	fe842783	;
assign	mem[11'd51]	=	32'h	00f707b3	;
assign	mem[11'd52]	=	32'h	0007c783	;
assign	mem[11'd53]	=	32'h	fe744703	;
assign	mem[11'd54]	=	32'h	00f71e63	;
assign	mem[11'd55]	=	32'h	fdc42703	;
assign	mem[11'd56]	=	32'h	fec42783	;
assign	mem[11'd57]	=	32'h	00f707b3	;
assign	mem[11'd58]	=	32'h	00078023	;
assign	mem[11'd59]	=	32'h	fdc42783	;
assign	mem[11'd60]	=	32'h	0680006f	;
assign	mem[11'd61]	=	32'h	fe842783	;
assign	mem[11'd62]	=	32'h	00178793	;
assign	mem[11'd63]	=	32'h	fef42423	;
assign	mem[11'd64]	=	32'h	fd442703	;
assign	mem[11'd65]	=	32'h	fe842783	;
assign	mem[11'd66]	=	32'h	00f707b3	;
assign	mem[11'd67]	=	32'h	0007c783	;
assign	mem[11'd68]	=	32'h	fa079ae3	;
assign	mem[11'd69]	=	32'h	fdc42703	;
assign	mem[11'd70]	=	32'h	fec42783	;
assign	mem[11'd71]	=	32'h	00f707b3	;
assign	mem[11'd72]	=	32'h	fe744703	;
assign	mem[11'd73]	=	32'h	00e78023	;
assign	mem[11'd74]	=	32'h	fec42783	;
assign	mem[11'd75]	=	32'h	00178793	;
assign	mem[11'd76]	=	32'h	fef42623	;
assign	mem[11'd77]	=	32'h	fec42703	;
assign	mem[11'd78]	=	32'h	fd842783	;
assign	mem[11'd79]	=	32'h	f6f76ae3	;
assign	mem[11'd80]	=	32'h	fd842783	;
assign	mem[11'd81]	=	32'h	fff78793	;
assign	mem[11'd82]	=	32'h	fdc42703	;
assign	mem[11'd83]	=	32'h	00f707b3	;
assign	mem[11'd84]	=	32'h	00078023	;
assign	mem[11'd85]	=	32'h	fdc42783	;
assign	mem[11'd86]	=	32'h	00078513	;
assign	mem[11'd87]	=	32'h	02c12083	;
assign	mem[11'd88]	=	32'h	02812403	;
assign	mem[11'd89]	=	32'h	03010113	;
assign	mem[11'd90]	=	32'h	00008067	;
assign	mem[11'd91]	=	32'h	fc010113	;
assign	mem[11'd92]	=	32'h	02112e23	;
assign	mem[11'd93]	=	32'h	02812c23	;
assign	mem[11'd94]	=	32'h	04010413	;
assign	mem[11'd95]	=	32'h	fca42623	;
assign	mem[11'd96]	=	32'h	fcb42423	;
assign	mem[11'd97]	=	32'h	fe042623	;
assign	mem[11'd98]	=	32'h	04c0006f	;
assign	mem[11'd99]	=	32'h	fd840793	;
assign	mem[11'd100]	=	32'h	00800593	;
assign	mem[11'd101]	=	32'h	00078513	;
assign	mem[11'd102]	=	32'h	e75ff0ef	;
assign	mem[11'd103]	=	32'h	fea42423	;
assign	mem[11'd104]	=	32'h	fec42783	;
assign	mem[11'd105]	=	32'h	00279713	;
assign	mem[11'd106]	=	32'h	fcc42783	;
assign	mem[11'd107]	=	32'h	00f707b3	;
assign	mem[11'd108]	=	32'h	fef42223	;
assign	mem[11'd109]	=	32'h	fe842503	;
assign	mem[11'd110]	=	32'h	0b9000ef	;
assign	mem[11'd111]	=	32'h	00050713	;
assign	mem[11'd112]	=	32'h	fe442783	;
assign	mem[11'd113]	=	32'h	00e7a023	;
assign	mem[11'd114]	=	32'h	fec42783	;
assign	mem[11'd115]	=	32'h	00178793	;
assign	mem[11'd116]	=	32'h	fef42623	;
assign	mem[11'd117]	=	32'h	fec42783	;
assign	mem[11'd118]	=	32'h	00279793	;
assign	mem[11'd119]	=	32'h	fc842703	;
assign	mem[11'd120]	=	32'h	fae7e6e3	;
assign	mem[11'd121]	=	32'h	00000013	;
assign	mem[11'd122]	=	32'h	03c12083	;
assign	mem[11'd123]	=	32'h	03812403	;
assign	mem[11'd124]	=	32'h	04010113	;
assign	mem[11'd125]	=	32'h	00008067	;
assign	mem[11'd126]	=	32'h	f4010113	;
assign	mem[11'd127]	=	32'h	0a112e23	;
assign	mem[11'd128]	=	32'h	0a812c23	;
assign	mem[11'd129]	=	32'h	0c010413	;
assign	mem[11'd130]	=	32'h	00001517	;
assign	mem[11'd131]	=	32'h	ea050513	;
assign	mem[11'd132]	=	32'h	5bd000ef	;
assign	mem[11'd133]	=	32'h	00001517	;
assign	mem[11'd134]	=	32'h	e9850513	;
assign	mem[11'd135]	=	32'h	5b1000ef	;
assign	mem[11'd136]	=	32'h	f4840793	;
assign	mem[11'd137]	=	32'h	00001617	;
assign	mem[11'd138]	=	32'h	e9060613	;
assign	mem[11'd139]	=	32'h	08000593	;
assign	mem[11'd140]	=	32'h	00078513	;
assign	mem[11'd141]	=	32'h	e59ff0ef	;
assign	mem[11'd142]	=	32'h	fea42623	;
assign	mem[11'd143]	=	32'h	00001597	;
assign	mem[11'd144]	=	32'h	e7c58593	;
assign	mem[11'd145]	=	32'h	fec42503	;
assign	mem[11'd146]	=	32'h	471000ef	;
assign	mem[11'd147]	=	32'h	00050793	;
assign	mem[11'd148]	=	32'h	06079263	;
assign	mem[11'd149]	=	32'h	f4840793	;
assign	mem[11'd150]	=	32'h	00001617	;
assign	mem[11'd151]	=	32'h	e5c60613	;
assign	mem[11'd152]	=	32'h	08000593	;
assign	mem[11'd153]	=	32'h	00078513	;
assign	mem[11'd154]	=	32'h	e25ff0ef	;
assign	mem[11'd155]	=	32'h	00050793	;
assign	mem[11'd156]	=	32'h	00078513	;
assign	mem[11'd157]	=	32'h	7fc000ef	;
assign	mem[11'd158]	=	32'h	fea42423	;
assign	mem[11'd159]	=	32'h	f4840793	;
assign	mem[11'd160]	=	32'h	00001617	;
assign	mem[11'd161]	=	32'h	e3460613	;
assign	mem[11'd162]	=	32'h	08000593	;
assign	mem[11'd163]	=	32'h	00078513	;
assign	mem[11'd164]	=	32'h	dfdff0ef	;
assign	mem[11'd165]	=	32'h	00050793	;
assign	mem[11'd166]	=	32'h	00078513	;
assign	mem[11'd167]	=	32'h	408000ef	;
assign	mem[11'd168]	=	32'h	fea42223	;
assign	mem[11'd169]	=	32'h	fe442583	;
assign	mem[11'd170]	=	32'h	fe842503	;
assign	mem[11'd171]	=	32'h	ec1ff0ef	;
assign	mem[11'd172]	=	32'h	f65ff06f	;
assign	mem[11'd173]	=	32'h	00001597	;
assign	mem[11'd174]	=	32'h	e0c58593	;
assign	mem[11'd175]	=	32'h	fec42503	;
assign	mem[11'd176]	=	32'h	3f9000ef	;
assign	mem[11'd177]	=	32'h	00050793	;
assign	mem[11'd178]	=	32'h	04079063	;
assign	mem[11'd179]	=	32'h	f4840793	;
assign	mem[11'd180]	=	32'h	00001617	;
assign	mem[11'd181]	=	32'h	de460613	;
assign	mem[11'd182]	=	32'h	08000593	;
assign	mem[11'd183]	=	32'h	00078513	;
assign	mem[11'd184]	=	32'h	dadff0ef	;
assign	mem[11'd185]	=	32'h	00050793	;
assign	mem[11'd186]	=	32'h	00078513	;
assign	mem[11'd187]	=	32'h	784000ef	;
assign	mem[11'd188]	=	32'h	fea42023	;
assign	mem[11'd189]	=	32'h	fe042783	;
assign	mem[11'd190]	=	32'h	fcf42e23	;
assign	mem[11'd191]	=	32'h	fdc42783	;
assign	mem[11'd192]	=	32'h	000780e7	;
assign	mem[11'd193]	=	32'h	f11ff06f	;
assign	mem[11'd194]	=	32'h	00001597	;
assign	mem[11'd195]	=	32'h	dbc58593	;
assign	mem[11'd196]	=	32'h	fec42503	;
assign	mem[11'd197]	=	32'h	3a5000ef	;
assign	mem[11'd198]	=	32'h	00050793	;
assign	mem[11'd199]	=	32'h	06079663	;
assign	mem[11'd200]	=	32'h	f4840793	;
assign	mem[11'd201]	=	32'h	00001617	;
assign	mem[11'd202]	=	32'h	d9060613	;
assign	mem[11'd203]	=	32'h	08000593	;
assign	mem[11'd204]	=	32'h	00078513	;
assign	mem[11'd205]	=	32'h	d59ff0ef	;
assign	mem[11'd206]	=	32'h	00050793	;
assign	mem[11'd207]	=	32'h	00078513	;
assign	mem[11'd208]	=	32'h	730000ef	;
assign	mem[11'd209]	=	32'h	fca42c23	;
assign	mem[11'd210]	=	32'h	fd842783	;
assign	mem[11'd211]	=	32'h	fcf42a23	;
assign	mem[11'd212]	=	32'h	fd442783	;
assign	mem[11'd213]	=	32'h	0007a783	;
assign	mem[11'd214]	=	32'h	f4840713	;
assign	mem[11'd215]	=	32'h	08000613	;
assign	mem[11'd216]	=	32'h	00070593	;
assign	mem[11'd217]	=	32'h	00078513	;
assign	mem[11'd218]	=	32'h	259000ef	;
assign	mem[11'd219]	=	32'h	00050793	;
assign	mem[11'd220]	=	32'h	00078513	;
assign	mem[11'd221]	=	32'h	459000ef	;
assign	mem[11'd222]	=	32'h	00001517	;
assign	mem[11'd223]	=	32'h	d3050513	;
assign	mem[11'd224]	=	32'h	44d000ef	;
assign	mem[11'd225]	=	32'h	e91ff06f	;
assign	mem[11'd226]	=	32'h	00001597	;
assign	mem[11'd227]	=	32'h	d4058593	;
assign	mem[11'd228]	=	32'h	fec42503	;
assign	mem[11'd229]	=	32'h	325000ef	;
assign	mem[11'd230]	=	32'h	00050793	;
assign	mem[11'd231]	=	32'h	06079663	;
assign	mem[11'd232]	=	32'h	f4840793	;
assign	mem[11'd233]	=	32'h	00001617	;
assign	mem[11'd234]	=	32'h	d1060613	;
assign	mem[11'd235]	=	32'h	08000593	;
assign	mem[11'd236]	=	32'h	00078513	;
assign	mem[11'd237]	=	32'h	cd9ff0ef	;
assign	mem[11'd238]	=	32'h	00050793	;
assign	mem[11'd239]	=	32'h	00078513	;
assign	mem[11'd240]	=	32'h	6b0000ef	;
assign	mem[11'd241]	=	32'h	fca42823	;
assign	mem[11'd242]	=	32'h	f4840793	;
assign	mem[11'd243]	=	32'h	00001617	;
assign	mem[11'd244]	=	32'h	ce860613	;
assign	mem[11'd245]	=	32'h	08000593	;
assign	mem[11'd246]	=	32'h	00078513	;
assign	mem[11'd247]	=	32'h	cb1ff0ef	;
assign	mem[11'd248]	=	32'h	00050793	;
assign	mem[11'd249]	=	32'h	00078513	;
assign	mem[11'd250]	=	32'h	688000ef	;
assign	mem[11'd251]	=	32'h	fca42623	;
assign	mem[11'd252]	=	32'h	fcc42783	;
assign	mem[11'd253]	=	32'h	fcf42423	;
assign	mem[11'd254]	=	32'h	fc842783	;
assign	mem[11'd255]	=	32'h	fd042703	;
assign	mem[11'd256]	=	32'h	00e7a023	;
assign	mem[11'd257]	=	32'h	e11ff06f	;
assign	mem[11'd258]	=	32'h	00001517	;
assign	mem[11'd259]	=	32'h	cc450513	;
assign	mem[11'd260]	=	32'h	3bd000ef	;
assign	mem[11'd261]	=	32'h	fec42503	;
assign	mem[11'd262]	=	32'h	3b5000ef	;
assign	mem[11'd263]	=	32'h	00001517	;
assign	mem[11'd264]	=	32'h	cbc50513	;
assign	mem[11'd265]	=	32'h	3a9000ef	;
assign	mem[11'd266]	=	32'h	dedff06f	;
assign	mem[11'd267]	=	32'h	fd010113	;
assign	mem[11'd268]	=	32'h	02812623	;
assign	mem[11'd269]	=	32'h	03010413	;
assign	mem[11'd270]	=	32'h	fca42e23	;
assign	mem[11'd271]	=	32'h	00058793	;
assign	mem[11'd272]	=	32'h	fcc42a23	;
assign	mem[11'd273]	=	32'h	fcf40da3	;
assign	mem[11'd274]	=	32'h	fe042623	;
assign	mem[11'd275]	=	32'h	0240006f	;
assign	mem[11'd276]	=	32'h	fdc42703	;
assign	mem[11'd277]	=	32'h	fec42783	;
assign	mem[11'd278]	=	32'h	00f707b3	;
assign	mem[11'd279]	=	32'h	fdb44703	;
assign	mem[11'd280]	=	32'h	00e78023	;
assign	mem[11'd281]	=	32'h	fec42783	;
assign	mem[11'd282]	=	32'h	00178793	;
assign	mem[11'd283]	=	32'h	fef42623	;
assign	mem[11'd284]	=	32'h	fec42703	;
assign	mem[11'd285]	=	32'h	fd442783	;
assign	mem[11'd286]	=	32'h	fcf76ce3	;
assign	mem[11'd287]	=	32'h	fdc42783	;
assign	mem[11'd288]	=	32'h	00078513	;
assign	mem[11'd289]	=	32'h	02c12403	;
assign	mem[11'd290]	=	32'h	03010113	;
assign	mem[11'd291]	=	32'h	00008067	;
assign	mem[11'd292]	=	32'h	fd010113	;
assign	mem[11'd293]	=	32'h	02812623	;
assign	mem[11'd294]	=	32'h	03010413	;
assign	mem[11'd295]	=	32'h	fca42e23	;
assign	mem[11'd296]	=	32'h	00058793	;
assign	mem[11'd297]	=	32'h	fcc42a23	;
assign	mem[11'd298]	=	32'h	fcf40da3	;
assign	mem[11'd299]	=	32'h	fe042623	;
assign	mem[11'd300]	=	32'h	0240006f	;
assign	mem[11'd301]	=	32'h	fdc42703	;
assign	mem[11'd302]	=	32'h	fec42783	;
assign	mem[11'd303]	=	32'h	00f707b3	;
assign	mem[11'd304]	=	32'h	fdb44703	;
assign	mem[11'd305]	=	32'h	00e78023	;
assign	mem[11'd306]	=	32'h	fec42783	;
assign	mem[11'd307]	=	32'h	00178793	;
assign	mem[11'd308]	=	32'h	fef42623	;
assign	mem[11'd309]	=	32'h	fec42703	;
assign	mem[11'd310]	=	32'h	fd442783	;
assign	mem[11'd311]	=	32'h	fcf76ce3	;
assign	mem[11'd312]	=	32'h	fdc42783	;
assign	mem[11'd313]	=	32'h	00078513	;
assign	mem[11'd314]	=	32'h	02c12403	;
assign	mem[11'd315]	=	32'h	03010113	;
assign	mem[11'd316]	=	32'h	00008067	;
assign	mem[11'd317]	=	32'h	fd010113	;
assign	mem[11'd318]	=	32'h	02812623	;
assign	mem[11'd319]	=	32'h	03010413	;
assign	mem[11'd320]	=	32'h	fca42e23	;
assign	mem[11'd321]	=	32'h	fe0407a3	;
assign	mem[11'd322]	=	32'h	fe042423	;
assign	mem[11'd323]	=	32'h	0800006f	;
assign	mem[11'd324]	=	32'h	fdc42703	;
assign	mem[11'd325]	=	32'h	fe842783	;
assign	mem[11'd326]	=	32'h	00f707b3	;
assign	mem[11'd327]	=	32'h	0007c703	;
assign	mem[11'd328]	=	32'h	02f00793	;
assign	mem[11'd329]	=	32'h	04e7fe63	;
assign	mem[11'd330]	=	32'h	fdc42703	;
assign	mem[11'd331]	=	32'h	fe842783	;
assign	mem[11'd332]	=	32'h	00f707b3	;
assign	mem[11'd333]	=	32'h	0007c703	;
assign	mem[11'd334]	=	32'h	03900793	;
assign	mem[11'd335]	=	32'h	04e7e263	;
assign	mem[11'd336]	=	32'h	fef44783	;
assign	mem[11'd337]	=	32'h	00379793	;
assign	mem[11'd338]	=	32'h	0ff7f713	;
assign	mem[11'd339]	=	32'h	fef44783	;
assign	mem[11'd340]	=	32'h	00179793	;
assign	mem[11'd341]	=	32'h	0ff7f793	;
assign	mem[11'd342]	=	32'h	00f707b3	;
assign	mem[11'd343]	=	32'h	0ff7f713	;
assign	mem[11'd344]	=	32'h	fdc42683	;
assign	mem[11'd345]	=	32'h	fe842783	;
assign	mem[11'd346]	=	32'h	00f687b3	;
assign	mem[11'd347]	=	32'h	0007c783	;
assign	mem[11'd348]	=	32'h	00f707b3	;
assign	mem[11'd349]	=	32'h	0ff7f793	;
assign	mem[11'd350]	=	32'h	fd078793	;
assign	mem[11'd351]	=	32'h	fef407a3	;
assign	mem[11'd352]	=	32'h	fe842783	;
assign	mem[11'd353]	=	32'h	00178793	;
assign	mem[11'd354]	=	32'h	fef42423	;
assign	mem[11'd355]	=	32'h	fe842703	;
assign	mem[11'd356]	=	32'h	00200793	;
assign	mem[11'd357]	=	32'h	00e7ec63	;
assign	mem[11'd358]	=	32'h	fdc42703	;
assign	mem[11'd359]	=	32'h	fe842783	;
assign	mem[11'd360]	=	32'h	00f707b3	;
assign	mem[11'd361]	=	32'h	0007c783	;
assign	mem[11'd362]	=	32'h	f60794e3	;
assign	mem[11'd363]	=	32'h	fef44783	;
assign	mem[11'd364]	=	32'h	00078513	;
assign	mem[11'd365]	=	32'h	02c12403	;
assign	mem[11'd366]	=	32'h	03010113	;
assign	mem[11'd367]	=	32'h	00008067	;
assign	mem[11'd368]	=	32'h	fd010113	;
assign	mem[11'd369]	=	32'h	02812623	;
assign	mem[11'd370]	=	32'h	03010413	;
assign	mem[11'd371]	=	32'h	fca42e23	;
assign	mem[11'd372]	=	32'h	fe041723	;
assign	mem[11'd373]	=	32'h	fe042423	;
assign	mem[11'd374]	=	32'h	0980006f	;
assign	mem[11'd375]	=	32'h	fdc42703	;
assign	mem[11'd376]	=	32'h	fe842783	;
assign	mem[11'd377]	=	32'h	00f707b3	;
assign	mem[11'd378]	=	32'h	0007c703	;
assign	mem[11'd379]	=	32'h	02f00793	;
assign	mem[11'd380]	=	32'h	06e7fa63	;
assign	mem[11'd381]	=	32'h	fdc42703	;
assign	mem[11'd382]	=	32'h	fe842783	;
assign	mem[11'd383]	=	32'h	00f707b3	;
assign	mem[11'd384]	=	32'h	0007c703	;
assign	mem[11'd385]	=	32'h	03900793	;
assign	mem[11'd386]	=	32'h	04e7ee63	;
assign	mem[11'd387]	=	32'h	fee45783	;
assign	mem[11'd388]	=	32'h	00379793	;
assign	mem[11'd389]	=	32'h	01079713	;
assign	mem[11'd390]	=	32'h	01075713	;
assign	mem[11'd391]	=	32'h	fee45783	;
assign	mem[11'd392]	=	32'h	00179793	;
assign	mem[11'd393]	=	32'h	01079793	;
assign	mem[11'd394]	=	32'h	0107d793	;
assign	mem[11'd395]	=	32'h	00f707b3	;
assign	mem[11'd396]	=	32'h	01079713	;
assign	mem[11'd397]	=	32'h	01075713	;
assign	mem[11'd398]	=	32'h	fdc42683	;
assign	mem[11'd399]	=	32'h	fe842783	;
assign	mem[11'd400]	=	32'h	00f687b3	;
assign	mem[11'd401]	=	32'h	0007c783	;
assign	mem[11'd402]	=	32'h	01079793	;
assign	mem[11'd403]	=	32'h	0107d793	;
assign	mem[11'd404]	=	32'h	00f707b3	;
assign	mem[11'd405]	=	32'h	01079793	;
assign	mem[11'd406]	=	32'h	0107d793	;
assign	mem[11'd407]	=	32'h	fd078793	;
assign	mem[11'd408]	=	32'h	fef41723	;
assign	mem[11'd409]	=	32'h	fe842783	;
assign	mem[11'd410]	=	32'h	00178793	;
assign	mem[11'd411]	=	32'h	fef42423	;
assign	mem[11'd412]	=	32'h	fe842703	;
assign	mem[11'd413]	=	32'h	00400793	;
assign	mem[11'd414]	=	32'h	00e7ec63	;
assign	mem[11'd415]	=	32'h	fdc42703	;
assign	mem[11'd416]	=	32'h	fe842783	;
assign	mem[11'd417]	=	32'h	00f707b3	;
assign	mem[11'd418]	=	32'h	0007c783	;
assign	mem[11'd419]	=	32'h	f40798e3	;
assign	mem[11'd420]	=	32'h	fee45783	;
assign	mem[11'd421]	=	32'h	00078513	;
assign	mem[11'd422]	=	32'h	02c12403	;
assign	mem[11'd423]	=	32'h	03010113	;
assign	mem[11'd424]	=	32'h	00008067	;
assign	mem[11'd425]	=	32'h	fd010113	;
assign	mem[11'd426]	=	32'h	02812623	;
assign	mem[11'd427]	=	32'h	03010413	;
assign	mem[11'd428]	=	32'h	fca42e23	;
assign	mem[11'd429]	=	32'h	fe042623	;
assign	mem[11'd430]	=	32'h	fe042423	;
assign	mem[11'd431]	=	32'h	0700006f	;
assign	mem[11'd432]	=	32'h	fdc42703	;
assign	mem[11'd433]	=	32'h	fe842783	;
assign	mem[11'd434]	=	32'h	00f707b3	;
assign	mem[11'd435]	=	32'h	0007c703	;
assign	mem[11'd436]	=	32'h	02f00793	;
assign	mem[11'd437]	=	32'h	04e7f663	;
assign	mem[11'd438]	=	32'h	fdc42703	;
assign	mem[11'd439]	=	32'h	fe842783	;
assign	mem[11'd440]	=	32'h	00f707b3	;
assign	mem[11'd441]	=	32'h	0007c703	;
assign	mem[11'd442]	=	32'h	03900793	;
assign	mem[11'd443]	=	32'h	02e7ea63	;
assign	mem[11'd444]	=	32'h	fec42783	;
assign	mem[11'd445]	=	32'h	00379713	;
assign	mem[11'd446]	=	32'h	fec42783	;
assign	mem[11'd447]	=	32'h	00179793	;
assign	mem[11'd448]	=	32'h	00f707b3	;
assign	mem[11'd449]	=	32'h	fdc42683	;
assign	mem[11'd450]	=	32'h	fe842703	;
assign	mem[11'd451]	=	32'h	00e68733	;
assign	mem[11'd452]	=	32'h	00074703	;
assign	mem[11'd453]	=	32'h	00e787b3	;
assign	mem[11'd454]	=	32'h	fd078793	;
assign	mem[11'd455]	=	32'h	fef42623	;
assign	mem[11'd456]	=	32'h	fe842783	;
assign	mem[11'd457]	=	32'h	00178793	;
assign	mem[11'd458]	=	32'h	fef42423	;
assign	mem[11'd459]	=	32'h	fe842703	;
assign	mem[11'd460]	=	32'h	00800793	;
assign	mem[11'd461]	=	32'h	00e7ec63	;
assign	mem[11'd462]	=	32'h	fdc42703	;
assign	mem[11'd463]	=	32'h	fe842783	;
assign	mem[11'd464]	=	32'h	00f707b3	;
assign	mem[11'd465]	=	32'h	0007c783	;
assign	mem[11'd466]	=	32'h	f6079ce3	;
assign	mem[11'd467]	=	32'h	fec42783	;
assign	mem[11'd468]	=	32'h	00078513	;
assign	mem[11'd469]	=	32'h	02c12403	;
assign	mem[11'd470]	=	32'h	03010113	;
assign	mem[11'd471]	=	32'h	00008067	;
assign	mem[11'd472]	=	32'h	fd010113	;
assign	mem[11'd473]	=	32'h	02812623	;
assign	mem[11'd474]	=	32'h	03010413	;
assign	mem[11'd475]	=	32'h	fca42e23	;
assign	mem[11'd476]	=	32'h	fe0407a3	;
assign	mem[11'd477]	=	32'h	fe040723	;
assign	mem[11'd478]	=	32'h	1240006f	;
assign	mem[11'd479]	=	32'h	fee44783	;
assign	mem[11'd480]	=	32'h	fdc42703	;
assign	mem[11'd481]	=	32'h	00f707b3	;
assign	mem[11'd482]	=	32'h	0007c703	;
assign	mem[11'd483]	=	32'h	02f00793	;
assign	mem[11'd484]	=	32'h	04e7f463	;
assign	mem[11'd485]	=	32'h	fee44783	;
assign	mem[11'd486]	=	32'h	fdc42703	;
assign	mem[11'd487]	=	32'h	00f707b3	;
assign	mem[11'd488]	=	32'h	0007c703	;
assign	mem[11'd489]	=	32'h	03900793	;
assign	mem[11'd490]	=	32'h	02e7e863	;
assign	mem[11'd491]	=	32'h	fef44783	;
assign	mem[11'd492]	=	32'h	00479793	;
assign	mem[11'd493]	=	32'h	0ff7f713	;
assign	mem[11'd494]	=	32'h	fee44783	;
assign	mem[11'd495]	=	32'h	fdc42683	;
assign	mem[11'd496]	=	32'h	00f687b3	;
assign	mem[11'd497]	=	32'h	0007c783	;
assign	mem[11'd498]	=	32'h	00f707b3	;
assign	mem[11'd499]	=	32'h	0ff7f793	;
assign	mem[11'd500]	=	32'h	fd078793	;
assign	mem[11'd501]	=	32'h	fef407a3	;
assign	mem[11'd502]	=	32'h	fee44783	;
assign	mem[11'd503]	=	32'h	fdc42703	;
assign	mem[11'd504]	=	32'h	00f707b3	;
assign	mem[11'd505]	=	32'h	0007c703	;
assign	mem[11'd506]	=	32'h	06000793	;
assign	mem[11'd507]	=	32'h	04e7f463	;
assign	mem[11'd508]	=	32'h	fee44783	;
assign	mem[11'd509]	=	32'h	fdc42703	;
assign	mem[11'd510]	=	32'h	00f707b3	;
assign	mem[11'd511]	=	32'h	0007c703	;
assign	mem[11'd512]	=	32'h	06600793	;
assign	mem[11'd513]	=	32'h	02e7e863	;
assign	mem[11'd514]	=	32'h	fef44783	;
assign	mem[11'd515]	=	32'h	00479793	;
assign	mem[11'd516]	=	32'h	0ff7f713	;
assign	mem[11'd517]	=	32'h	fee44783	;
assign	mem[11'd518]	=	32'h	fdc42683	;
assign	mem[11'd519]	=	32'h	00f687b3	;
assign	mem[11'd520]	=	32'h	0007c783	;
assign	mem[11'd521]	=	32'h	00f707b3	;
assign	mem[11'd522]	=	32'h	0ff7f793	;
assign	mem[11'd523]	=	32'h	fa978793	;
assign	mem[11'd524]	=	32'h	fef407a3	;
assign	mem[11'd525]	=	32'h	fee44783	;
assign	mem[11'd526]	=	32'h	fdc42703	;
assign	mem[11'd527]	=	32'h	00f707b3	;
assign	mem[11'd528]	=	32'h	0007c703	;
assign	mem[11'd529]	=	32'h	04000793	;
assign	mem[11'd530]	=	32'h	04e7f463	;
assign	mem[11'd531]	=	32'h	fee44783	;
assign	mem[11'd532]	=	32'h	fdc42703	;
assign	mem[11'd533]	=	32'h	00f707b3	;
assign	mem[11'd534]	=	32'h	0007c703	;
assign	mem[11'd535]	=	32'h	04600793	;
assign	mem[11'd536]	=	32'h	02e7e863	;
assign	mem[11'd537]	=	32'h	fef44783	;
assign	mem[11'd538]	=	32'h	00479793	;
assign	mem[11'd539]	=	32'h	0ff7f713	;
assign	mem[11'd540]	=	32'h	fee44783	;
assign	mem[11'd541]	=	32'h	fdc42683	;
assign	mem[11'd542]	=	32'h	00f687b3	;
assign	mem[11'd543]	=	32'h	0007c783	;
assign	mem[11'd544]	=	32'h	00f707b3	;
assign	mem[11'd545]	=	32'h	0ff7f793	;
assign	mem[11'd546]	=	32'h	fc978793	;
assign	mem[11'd547]	=	32'h	fef407a3	;
assign	mem[11'd548]	=	32'h	fee44783	;
assign	mem[11'd549]	=	32'h	00178793	;
assign	mem[11'd550]	=	32'h	fef40723	;
assign	mem[11'd551]	=	32'h	fee44703	;
assign	mem[11'd552]	=	32'h	00100793	;
assign	mem[11'd553]	=	32'h	00e7ec63	;
assign	mem[11'd554]	=	32'h	fee44783	;
assign	mem[11'd555]	=	32'h	fdc42703	;
assign	mem[11'd556]	=	32'h	00f707b3	;
assign	mem[11'd557]	=	32'h	0007c783	;
assign	mem[11'd558]	=	32'h	ec0792e3	;
assign	mem[11'd559]	=	32'h	fef44783	;
assign	mem[11'd560]	=	32'h	00078513	;
assign	mem[11'd561]	=	32'h	02c12403	;
assign	mem[11'd562]	=	32'h	03010113	;
assign	mem[11'd563]	=	32'h	00008067	;
assign	mem[11'd564]	=	32'h	fd010113	;
assign	mem[11'd565]	=	32'h	02812623	;
assign	mem[11'd566]	=	32'h	03010413	;
assign	mem[11'd567]	=	32'h	fca42e23	;
assign	mem[11'd568]	=	32'h	fe041723	;
assign	mem[11'd569]	=	32'h	fe041623	;
assign	mem[11'd570]	=	32'h	1540006f	;
assign	mem[11'd571]	=	32'h	fec45783	;
assign	mem[11'd572]	=	32'h	fdc42703	;
assign	mem[11'd573]	=	32'h	00f707b3	;
assign	mem[11'd574]	=	32'h	0007c703	;
assign	mem[11'd575]	=	32'h	02f00793	;
assign	mem[11'd576]	=	32'h	04e7fc63	;
assign	mem[11'd577]	=	32'h	fec45783	;
assign	mem[11'd578]	=	32'h	fdc42703	;
assign	mem[11'd579]	=	32'h	00f707b3	;
assign	mem[11'd580]	=	32'h	0007c703	;
assign	mem[11'd581]	=	32'h	03900793	;
assign	mem[11'd582]	=	32'h	04e7e063	;
assign	mem[11'd583]	=	32'h	fee45783	;
assign	mem[11'd584]	=	32'h	00479793	;
assign	mem[11'd585]	=	32'h	01079713	;
assign	mem[11'd586]	=	32'h	01075713	;
assign	mem[11'd587]	=	32'h	fec45783	;
assign	mem[11'd588]	=	32'h	fdc42683	;
assign	mem[11'd589]	=	32'h	00f687b3	;
assign	mem[11'd590]	=	32'h	0007c783	;
assign	mem[11'd591]	=	32'h	01079793	;
assign	mem[11'd592]	=	32'h	0107d793	;
assign	mem[11'd593]	=	32'h	00f707b3	;
assign	mem[11'd594]	=	32'h	01079793	;
assign	mem[11'd595]	=	32'h	0107d793	;
assign	mem[11'd596]	=	32'h	fd078793	;
assign	mem[11'd597]	=	32'h	fef41723	;
assign	mem[11'd598]	=	32'h	fec45783	;
assign	mem[11'd599]	=	32'h	fdc42703	;
assign	mem[11'd600]	=	32'h	00f707b3	;
assign	mem[11'd601]	=	32'h	0007c703	;
assign	mem[11'd602]	=	32'h	06000793	;
assign	mem[11'd603]	=	32'h	04e7fc63	;
assign	mem[11'd604]	=	32'h	fec45783	;
assign	mem[11'd605]	=	32'h	fdc42703	;
assign	mem[11'd606]	=	32'h	00f707b3	;
assign	mem[11'd607]	=	32'h	0007c703	;
assign	mem[11'd608]	=	32'h	06600793	;
assign	mem[11'd609]	=	32'h	04e7e063	;
assign	mem[11'd610]	=	32'h	fee45783	;
assign	mem[11'd611]	=	32'h	00479793	;
assign	mem[11'd612]	=	32'h	01079713	;
assign	mem[11'd613]	=	32'h	01075713	;
assign	mem[11'd614]	=	32'h	fec45783	;
assign	mem[11'd615]	=	32'h	fdc42683	;
assign	mem[11'd616]	=	32'h	00f687b3	;
assign	mem[11'd617]	=	32'h	0007c783	;
assign	mem[11'd618]	=	32'h	01079793	;
assign	mem[11'd619]	=	32'h	0107d793	;
assign	mem[11'd620]	=	32'h	00f707b3	;
assign	mem[11'd621]	=	32'h	01079793	;
assign	mem[11'd622]	=	32'h	0107d793	;
assign	mem[11'd623]	=	32'h	fa978793	;
assign	mem[11'd624]	=	32'h	fef41723	;
assign	mem[11'd625]	=	32'h	fec45783	;
assign	mem[11'd626]	=	32'h	fdc42703	;
assign	mem[11'd627]	=	32'h	00f707b3	;
assign	mem[11'd628]	=	32'h	0007c703	;
assign	mem[11'd629]	=	32'h	04000793	;
assign	mem[11'd630]	=	32'h	04e7fc63	;
assign	mem[11'd631]	=	32'h	fec45783	;
assign	mem[11'd632]	=	32'h	fdc42703	;
assign	mem[11'd633]	=	32'h	00f707b3	;
assign	mem[11'd634]	=	32'h	0007c703	;
assign	mem[11'd635]	=	32'h	04600793	;
assign	mem[11'd636]	=	32'h	04e7e063	;
assign	mem[11'd637]	=	32'h	fee45783	;
assign	mem[11'd638]	=	32'h	00479793	;
assign	mem[11'd639]	=	32'h	01079713	;
assign	mem[11'd640]	=	32'h	01075713	;
assign	mem[11'd641]	=	32'h	fec45783	;
assign	mem[11'd642]	=	32'h	fdc42683	;
assign	mem[11'd643]	=	32'h	00f687b3	;
assign	mem[11'd644]	=	32'h	0007c783	;
assign	mem[11'd645]	=	32'h	01079793	;
assign	mem[11'd646]	=	32'h	0107d793	;
assign	mem[11'd647]	=	32'h	00f707b3	;
assign	mem[11'd648]	=	32'h	01079793	;
assign	mem[11'd649]	=	32'h	0107d793	;
assign	mem[11'd650]	=	32'h	fc978793	;
assign	mem[11'd651]	=	32'h	fef41723	;
assign	mem[11'd652]	=	32'h	fec45783	;
assign	mem[11'd653]	=	32'h	00178793	;
assign	mem[11'd654]	=	32'h	fef41623	;
assign	mem[11'd655]	=	32'h	fec45703	;
assign	mem[11'd656]	=	32'h	00300793	;
assign	mem[11'd657]	=	32'h	00e7ec63	;
assign	mem[11'd658]	=	32'h	fec45783	;
assign	mem[11'd659]	=	32'h	fdc42703	;
assign	mem[11'd660]	=	32'h	00f707b3	;
assign	mem[11'd661]	=	32'h	0007c783	;
assign	mem[11'd662]	=	32'h	e8079ae3	;
assign	mem[11'd663]	=	32'h	fee45783	;
assign	mem[11'd664]	=	32'h	00078513	;
assign	mem[11'd665]	=	32'h	02c12403	;
assign	mem[11'd666]	=	32'h	03010113	;
assign	mem[11'd667]	=	32'h	00008067	;
assign	mem[11'd668]	=	32'h	fd010113	;
assign	mem[11'd669]	=	32'h	02812623	;
assign	mem[11'd670]	=	32'h	03010413	;
assign	mem[11'd671]	=	32'h	fca42e23	;
assign	mem[11'd672]	=	32'h	fe042623	;
assign	mem[11'd673]	=	32'h	fe042423	;
assign	mem[11'd674]	=	32'h	10c0006f	;
assign	mem[11'd675]	=	32'h	fdc42703	;
assign	mem[11'd676]	=	32'h	fe842783	;
assign	mem[11'd677]	=	32'h	00f707b3	;
assign	mem[11'd678]	=	32'h	0007c703	;
assign	mem[11'd679]	=	32'h	02f00793	;
assign	mem[11'd680]	=	32'h	04e7f063	;
assign	mem[11'd681]	=	32'h	fdc42703	;
assign	mem[11'd682]	=	32'h	fe842783	;
assign	mem[11'd683]	=	32'h	00f707b3	;
assign	mem[11'd684]	=	32'h	0007c703	;
assign	mem[11'd685]	=	32'h	03900793	;
assign	mem[11'd686]	=	32'h	02e7e463	;
assign	mem[11'd687]	=	32'h	fec42783	;
assign	mem[11'd688]	=	32'h	00479793	;
assign	mem[11'd689]	=	32'h	fdc42683	;
assign	mem[11'd690]	=	32'h	fe842703	;
assign	mem[11'd691]	=	32'h	00e68733	;
assign	mem[11'd692]	=	32'h	00074703	;
assign	mem[11'd693]	=	32'h	00e787b3	;
assign	mem[11'd694]	=	32'h	fd078793	;
assign	mem[11'd695]	=	32'h	fef42623	;
assign	mem[11'd696]	=	32'h	fdc42703	;
assign	mem[11'd697]	=	32'h	fe842783	;
assign	mem[11'd698]	=	32'h	00f707b3	;
assign	mem[11'd699]	=	32'h	0007c703	;
assign	mem[11'd700]	=	32'h	06000793	;
assign	mem[11'd701]	=	32'h	04e7f063	;
assign	mem[11'd702]	=	32'h	fdc42703	;
assign	mem[11'd703]	=	32'h	fe842783	;
assign	mem[11'd704]	=	32'h	00f707b3	;
assign	mem[11'd705]	=	32'h	0007c703	;
assign	mem[11'd706]	=	32'h	06600793	;
assign	mem[11'd707]	=	32'h	02e7e463	;
assign	mem[11'd708]	=	32'h	fec42783	;
assign	mem[11'd709]	=	32'h	00479793	;
assign	mem[11'd710]	=	32'h	fdc42683	;
assign	mem[11'd711]	=	32'h	fe842703	;
assign	mem[11'd712]	=	32'h	00e68733	;
assign	mem[11'd713]	=	32'h	00074703	;
assign	mem[11'd714]	=	32'h	00e787b3	;
assign	mem[11'd715]	=	32'h	fa978793	;
assign	mem[11'd716]	=	32'h	fef42623	;
assign	mem[11'd717]	=	32'h	fdc42703	;
assign	mem[11'd718]	=	32'h	fe842783	;
assign	mem[11'd719]	=	32'h	00f707b3	;
assign	mem[11'd720]	=	32'h	0007c703	;
assign	mem[11'd721]	=	32'h	04000793	;
assign	mem[11'd722]	=	32'h	04e7f063	;
assign	mem[11'd723]	=	32'h	fdc42703	;
assign	mem[11'd724]	=	32'h	fe842783	;
assign	mem[11'd725]	=	32'h	00f707b3	;
assign	mem[11'd726]	=	32'h	0007c703	;
assign	mem[11'd727]	=	32'h	04600793	;
assign	mem[11'd728]	=	32'h	02e7e463	;
assign	mem[11'd729]	=	32'h	fec42783	;
assign	mem[11'd730]	=	32'h	00479793	;
assign	mem[11'd731]	=	32'h	fdc42683	;
assign	mem[11'd732]	=	32'h	fe842703	;
assign	mem[11'd733]	=	32'h	00e68733	;
assign	mem[11'd734]	=	32'h	00074703	;
assign	mem[11'd735]	=	32'h	00e787b3	;
assign	mem[11'd736]	=	32'h	fc978793	;
assign	mem[11'd737]	=	32'h	fef42623	;
assign	mem[11'd738]	=	32'h	fe842783	;
assign	mem[11'd739]	=	32'h	00178793	;
assign	mem[11'd740]	=	32'h	fef42423	;
assign	mem[11'd741]	=	32'h	fe842703	;
assign	mem[11'd742]	=	32'h	00700793	;
assign	mem[11'd743]	=	32'h	00e7ec63	;
assign	mem[11'd744]	=	32'h	fdc42703	;
assign	mem[11'd745]	=	32'h	fe842783	;
assign	mem[11'd746]	=	32'h	00f707b3	;
assign	mem[11'd747]	=	32'h	0007c783	;
assign	mem[11'd748]	=	32'h	ec079ee3	;
assign	mem[11'd749]	=	32'h	fec42783	;
assign	mem[11'd750]	=	32'h	00078513	;
assign	mem[11'd751]	=	32'h	02c12403	;
assign	mem[11'd752]	=	32'h	03010113	;
assign	mem[11'd753]	=	32'h	00008067	;
assign	mem[11'd754]	=	32'h	fd010113	;
assign	mem[11'd755]	=	32'h	02812623	;
assign	mem[11'd756]	=	32'h	03010413	;
assign	mem[11'd757]	=	32'h	00050793	;
assign	mem[11'd758]	=	32'h	fcb42c23	;
assign	mem[11'd759]	=	32'h	fcc42a23	;
assign	mem[11'd760]	=	32'h	fcf40fa3	;
assign	mem[11'd761]	=	32'h	fe042623	;
assign	mem[11'd762]	=	32'h	00200793	;
assign	mem[11'd763]	=	32'h	fef42423	;
assign	mem[11'd764]	=	32'h	0940006f	;
assign	mem[11'd765]	=	32'h	fdf44703	;
assign	mem[11'd766]	=	32'h	fe842683	;
assign	mem[11'd767]	=	32'h	fec42783	;
assign	mem[11'd768]	=	32'h	40f687b3	;
assign	mem[11'd769]	=	32'h	fff78793	;
assign	mem[11'd770]	=	32'h	00279793	;
assign	mem[11'd771]	=	32'h	40f757b3	;
assign	mem[11'd772]	=	32'h	0ff7f793	;
assign	mem[11'd773]	=	32'h	00f7f793	;
assign	mem[11'd774]	=	32'h	fef403a3	;
assign	mem[11'd775]	=	32'h	fe744703	;
assign	mem[11'd776]	=	32'h	00900793	;
assign	mem[11'd777]	=	32'h	02e7e063	;
assign	mem[11'd778]	=	32'h	fd842703	;
assign	mem[11'd779]	=	32'h	fec42783	;
assign	mem[11'd780]	=	32'h	00f707b3	;
assign	mem[11'd781]	=	32'h	fe744703	;
assign	mem[11'd782]	=	32'h	03070713	;
assign	mem[11'd783]	=	32'h	0ff77713	;
assign	mem[11'd784]	=	32'h	00e78023	;
assign	mem[11'd785]	=	32'h	fe744703	;
assign	mem[11'd786]	=	32'h	00900793	;
assign	mem[11'd787]	=	32'h	02e7f663	;
assign	mem[11'd788]	=	32'h	fe744703	;
assign	mem[11'd789]	=	32'h	00f00793	;
assign	mem[11'd790]	=	32'h	02e7e063	;
assign	mem[11'd791]	=	32'h	fd842703	;
assign	mem[11'd792]	=	32'h	fec42783	;
assign	mem[11'd793]	=	32'h	00f707b3	;
assign	mem[11'd794]	=	32'h	fe744703	;
assign	mem[11'd795]	=	32'h	05770713	;
assign	mem[11'd796]	=	32'h	0ff77713	;
assign	mem[11'd797]	=	32'h	00e78023	;
assign	mem[11'd798]	=	32'h	fec42783	;
assign	mem[11'd799]	=	32'h	00178793	;
assign	mem[11'd800]	=	32'h	fef42623	;
assign	mem[11'd801]	=	32'h	fec42703	;
assign	mem[11'd802]	=	32'h	fe842783	;
assign	mem[11'd803]	=	32'h	00f77a63	;
assign	mem[11'd804]	=	32'h	fec42783	;
assign	mem[11'd805]	=	32'h	00178793	;
assign	mem[11'd806]	=	32'h	fd442703	;
assign	mem[11'd807]	=	32'h	f4e7ece3	;
assign	mem[11'd808]	=	32'h	fd842703	;
assign	mem[11'd809]	=	32'h	fec42783	;
assign	mem[11'd810]	=	32'h	00f707b3	;
assign	mem[11'd811]	=	32'h	00078023	;
assign	mem[11'd812]	=	32'h	fd842783	;
assign	mem[11'd813]	=	32'h	00078513	;
assign	mem[11'd814]	=	32'h	02c12403	;
assign	mem[11'd815]	=	32'h	03010113	;
assign	mem[11'd816]	=	32'h	00008067	;
assign	mem[11'd817]	=	32'h	fd010113	;
assign	mem[11'd818]	=	32'h	02812623	;
assign	mem[11'd819]	=	32'h	03010413	;
assign	mem[11'd820]	=	32'h	00050793	;
assign	mem[11'd821]	=	32'h	fcb42c23	;
assign	mem[11'd822]	=	32'h	fcc42a23	;
assign	mem[11'd823]	=	32'h	fcf41f23	;
assign	mem[11'd824]	=	32'h	fe042623	;
assign	mem[11'd825]	=	32'h	00400793	;
assign	mem[11'd826]	=	32'h	fef42423	;
assign	mem[11'd827]	=	32'h	0940006f	;
assign	mem[11'd828]	=	32'h	fde45703	;
assign	mem[11'd829]	=	32'h	fe842683	;
assign	mem[11'd830]	=	32'h	fec42783	;
assign	mem[11'd831]	=	32'h	40f687b3	;
assign	mem[11'd832]	=	32'h	fff78793	;
assign	mem[11'd833]	=	32'h	00279793	;
assign	mem[11'd834]	=	32'h	40f757b3	;
assign	mem[11'd835]	=	32'h	0ff7f793	;
assign	mem[11'd836]	=	32'h	00f7f793	;
assign	mem[11'd837]	=	32'h	fef403a3	;
assign	mem[11'd838]	=	32'h	fe744703	;
assign	mem[11'd839]	=	32'h	00900793	;
assign	mem[11'd840]	=	32'h	02e7e063	;
assign	mem[11'd841]	=	32'h	fd842703	;
assign	mem[11'd842]	=	32'h	fec42783	;
assign	mem[11'd843]	=	32'h	00f707b3	;
assign	mem[11'd844]	=	32'h	fe744703	;
assign	mem[11'd845]	=	32'h	03070713	;
assign	mem[11'd846]	=	32'h	0ff77713	;
assign	mem[11'd847]	=	32'h	00e78023	;
assign	mem[11'd848]	=	32'h	fe744703	;
assign	mem[11'd849]	=	32'h	00900793	;
assign	mem[11'd850]	=	32'h	02e7f663	;
assign	mem[11'd851]	=	32'h	fe744703	;
assign	mem[11'd852]	=	32'h	00f00793	;
assign	mem[11'd853]	=	32'h	02e7e063	;
assign	mem[11'd854]	=	32'h	fd842703	;
assign	mem[11'd855]	=	32'h	fec42783	;
assign	mem[11'd856]	=	32'h	00f707b3	;
assign	mem[11'd857]	=	32'h	fe744703	;
assign	mem[11'd858]	=	32'h	05770713	;
assign	mem[11'd859]	=	32'h	0ff77713	;
assign	mem[11'd860]	=	32'h	00e78023	;
assign	mem[11'd861]	=	32'h	fec42783	;
assign	mem[11'd862]	=	32'h	00178793	;
assign	mem[11'd863]	=	32'h	fef42623	;
assign	mem[11'd864]	=	32'h	fec42703	;
assign	mem[11'd865]	=	32'h	fe842783	;
assign	mem[11'd866]	=	32'h	00f77a63	;
assign	mem[11'd867]	=	32'h	fec42783	;
assign	mem[11'd868]	=	32'h	00178793	;
assign	mem[11'd869]	=	32'h	fd442703	;
assign	mem[11'd870]	=	32'h	f4e7ece3	;
assign	mem[11'd871]	=	32'h	fd842703	;
assign	mem[11'd872]	=	32'h	fec42783	;
assign	mem[11'd873]	=	32'h	00f707b3	;
assign	mem[11'd874]	=	32'h	00078023	;
assign	mem[11'd875]	=	32'h	fd842783	;
assign	mem[11'd876]	=	32'h	00078513	;
assign	mem[11'd877]	=	32'h	02c12403	;
assign	mem[11'd878]	=	32'h	03010113	;
assign	mem[11'd879]	=	32'h	00008067	;
assign	mem[11'd880]	=	32'h	fd010113	;
assign	mem[11'd881]	=	32'h	02812623	;
assign	mem[11'd882]	=	32'h	03010413	;
assign	mem[11'd883]	=	32'h	fca42e23	;
assign	mem[11'd884]	=	32'h	fcb42c23	;
assign	mem[11'd885]	=	32'h	fcc42a23	;
assign	mem[11'd886]	=	32'h	fe042623	;
assign	mem[11'd887]	=	32'h	00800793	;
assign	mem[11'd888]	=	32'h	fef42423	;
assign	mem[11'd889]	=	32'h	0940006f	;
assign	mem[11'd890]	=	32'h	fe842703	;
assign	mem[11'd891]	=	32'h	fec42783	;
assign	mem[11'd892]	=	32'h	40f707b3	;
assign	mem[11'd893]	=	32'h	fff78793	;
assign	mem[11'd894]	=	32'h	00279793	;
assign	mem[11'd895]	=	32'h	fdc42703	;
assign	mem[11'd896]	=	32'h	00f757b3	;
assign	mem[11'd897]	=	32'h	0ff7f793	;
assign	mem[11'd898]	=	32'h	00f7f793	;
assign	mem[11'd899]	=	32'h	fef403a3	;
assign	mem[11'd900]	=	32'h	fe744703	;
assign	mem[11'd901]	=	32'h	00900793	;
assign	mem[11'd902]	=	32'h	02e7e063	;
assign	mem[11'd903]	=	32'h	fd842703	;
assign	mem[11'd904]	=	32'h	fec42783	;
assign	mem[11'd905]	=	32'h	00f707b3	;
assign	mem[11'd906]	=	32'h	fe744703	;
assign	mem[11'd907]	=	32'h	03070713	;
assign	mem[11'd908]	=	32'h	0ff77713	;
assign	mem[11'd909]	=	32'h	00e78023	;
assign	mem[11'd910]	=	32'h	fe744703	;
assign	mem[11'd911]	=	32'h	00900793	;
assign	mem[11'd912]	=	32'h	02e7f663	;
assign	mem[11'd913]	=	32'h	fe744703	;
assign	mem[11'd914]	=	32'h	00f00793	;
assign	mem[11'd915]	=	32'h	02e7e063	;
assign	mem[11'd916]	=	32'h	fd842703	;
assign	mem[11'd917]	=	32'h	fec42783	;
assign	mem[11'd918]	=	32'h	00f707b3	;
assign	mem[11'd919]	=	32'h	fe744703	;
assign	mem[11'd920]	=	32'h	05770713	;
assign	mem[11'd921]	=	32'h	0ff77713	;
assign	mem[11'd922]	=	32'h	00e78023	;
assign	mem[11'd923]	=	32'h	fec42783	;
assign	mem[11'd924]	=	32'h	00178793	;
assign	mem[11'd925]	=	32'h	fef42623	;
assign	mem[11'd926]	=	32'h	fec42703	;
assign	mem[11'd927]	=	32'h	fe842783	;
assign	mem[11'd928]	=	32'h	00f77a63	;
assign	mem[11'd929]	=	32'h	fec42783	;
assign	mem[11'd930]	=	32'h	00178793	;
assign	mem[11'd931]	=	32'h	fd442703	;
assign	mem[11'd932]	=	32'h	f4e7ece3	;
assign	mem[11'd933]	=	32'h	fd842703	;
assign	mem[11'd934]	=	32'h	fec42783	;
assign	mem[11'd935]	=	32'h	00f707b3	;
assign	mem[11'd936]	=	32'h	00078023	;
assign	mem[11'd937]	=	32'h	fd842783	;
assign	mem[11'd938]	=	32'h	00078513	;
assign	mem[11'd939]	=	32'h	02c12403	;
assign	mem[11'd940]	=	32'h	03010113	;
assign	mem[11'd941]	=	32'h	00008067	;
assign	mem[11'd942]	=	32'h	fd010113	;
assign	mem[11'd943]	=	32'h	02812623	;
assign	mem[11'd944]	=	32'h	03010413	;
assign	mem[11'd945]	=	32'h	fca42e23	;
assign	mem[11'd946]	=	32'h	fcb42c23	;
assign	mem[11'd947]	=	32'h	fe042623	;
assign	mem[11'd948]	=	32'h	fdc42703	;
assign	mem[11'd949]	=	32'h	fec42783	;
assign	mem[11'd950]	=	32'h	00f707b3	;
assign	mem[11'd951]	=	32'h	0007c703	;
assign	mem[11'd952]	=	32'h	fd842683	;
assign	mem[11'd953]	=	32'h	fec42783	;
assign	mem[11'd954]	=	32'h	00f687b3	;
assign	mem[11'd955]	=	32'h	0007c783	;
assign	mem[11'd956]	=	32'h	00f70663	;
assign	mem[11'd957]	=	32'h	00100793	;
assign	mem[11'd958]	=	32'h	0300006f	;
assign	mem[11'd959]	=	32'h	fdc42703	;
assign	mem[11'd960]	=	32'h	fec42783	;
assign	mem[11'd961]	=	32'h	00f707b3	;
assign	mem[11'd962]	=	32'h	0007c783	;
assign	mem[11'd963]	=	32'h	00078a63	;
assign	mem[11'd964]	=	32'h	fec42783	;
assign	mem[11'd965]	=	32'h	00178793	;
assign	mem[11'd966]	=	32'h	fef42623	;
assign	mem[11'd967]	=	32'h	fb5ff06f	;
assign	mem[11'd968]	=	32'h	00000013	;
assign	mem[11'd969]	=	32'h	00000793	;
assign	mem[11'd970]	=	32'h	00078513	;
assign	mem[11'd971]	=	32'h	02c12403	;
assign	mem[11'd972]	=	32'h	03010113	;
assign	mem[11'd973]	=	32'h	00008067	;
assign	mem[11'd974]	=	32'h	fd010113	;
assign	mem[11'd975]	=	32'h	02812623	;
assign	mem[11'd976]	=	32'h	03010413	;
assign	mem[11'd977]	=	32'h	fca42e23	;
assign	mem[11'd978]	=	32'h	fe042623	;
assign	mem[11'd979]	=	32'h	0100006f	;
assign	mem[11'd980]	=	32'h	fec42783	;
assign	mem[11'd981]	=	32'h	00178793	;
assign	mem[11'd982]	=	32'h	fef42623	;
assign	mem[11'd983]	=	32'h	fdc42703	;
assign	mem[11'd984]	=	32'h	fec42783	;
assign	mem[11'd985]	=	32'h	00f707b3	;
assign	mem[11'd986]	=	32'h	0007c783	;
assign	mem[11'd987]	=	32'h	fe0792e3	;
assign	mem[11'd988]	=	32'h	fec42783	;
assign	mem[11'd989]	=	32'h	00078513	;
assign	mem[11'd990]	=	32'h	02c12403	;
assign	mem[11'd991]	=	32'h	03010113	;
assign	mem[11'd992]	=	32'h	00008067	;
assign	mem[11'd993]	=	32'h	fe010113	;
assign	mem[11'd994]	=	32'h	00812e23	;
assign	mem[11'd995]	=	32'h	02010413	;
assign	mem[11'd996]	=	32'h	00050793	;
assign	mem[11'd997]	=	32'h	fef407a3	;
assign	mem[11'd998]	=	32'h	00000013	;
assign	mem[11'd999]	=	32'h	800007b7	;
assign	mem[11'd1000]	=	32'h	0007a783	;
assign	mem[11'd1001]	=	32'h	0017f793	;
assign	mem[11'd1002]	=	32'h	fe078ae3	;
assign	mem[11'd1003]	=	32'h	800007b7	;
assign	mem[11'd1004]	=	32'h	00878793	;
assign	mem[11'd1005]	=	32'h	fef44703	;
assign	mem[11'd1006]	=	32'h	00e7a023	;
assign	mem[11'd1007]	=	32'h	00000013	;
assign	mem[11'd1008]	=	32'h	01c12403	;
assign	mem[11'd1009]	=	32'h	02010113	;
assign	mem[11'd1010]	=	32'h	00008067	;
assign	mem[11'd1011]	=	32'h	fd010113	;
assign	mem[11'd1012]	=	32'h	02112623	;
assign	mem[11'd1013]	=	32'h	02812423	;
assign	mem[11'd1014]	=	32'h	03010413	;
assign	mem[11'd1015]	=	32'h	fca42e23	;
assign	mem[11'd1016]	=	32'h	fe042623	;
assign	mem[11'd1017]	=	32'h	0280006f	;
assign	mem[11'd1018]	=	32'h	fec42783	;
assign	mem[11'd1019]	=	32'h	fdc42703	;
assign	mem[11'd1020]	=	32'h	00f707b3	;
assign	mem[11'd1021]	=	32'h	0007c783	;
assign	mem[11'd1022]	=	32'h	00078513	;
assign	mem[11'd1023]	=	32'h	f89ff0ef	;
assign	mem[11'd1024]	=	32'h	fec42783	;
assign	mem[11'd1025]	=	32'h	00178793	;
assign	mem[11'd1026]	=	32'h	fef42623	;
assign	mem[11'd1027]	=	32'h	fec42783	;
assign	mem[11'd1028]	=	32'h	fdc42703	;
assign	mem[11'd1029]	=	32'h	00f707b3	;
assign	mem[11'd1030]	=	32'h	0007c783	;
assign	mem[11'd1031]	=	32'h	fc0796e3	;
assign	mem[11'd1032]	=	32'h	00000013	;
assign	mem[11'd1033]	=	32'h	02c12083	;
assign	mem[11'd1034]	=	32'h	02812403	;
assign	mem[11'd1035]	=	32'h	03010113	;
assign	mem[11'd1036]	=	32'h	00008067	;
assign	mem[11'd1037]	=	32'h	fe010113	;
assign	mem[11'd1038]	=	32'h	00112e23	;
assign	mem[11'd1039]	=	32'h	00812c23	;
assign	mem[11'd1040]	=	32'h	02010413	;
assign	mem[11'd1041]	=	32'h	00000013	;
assign	mem[11'd1042]	=	32'h	800007b7	;
assign	mem[11'd1043]	=	32'h	0007a783	;
assign	mem[11'd1044]	=	32'h	0027f793	;
assign	mem[11'd1045]	=	32'h	fe078ae3	;
assign	mem[11'd1046]	=	32'h	800007b7	;
assign	mem[11'd1047]	=	32'h	00478793	;
assign	mem[11'd1048]	=	32'h	0007a783	;
assign	mem[11'd1049]	=	32'h	fef407a3	;
assign	mem[11'd1050]	=	32'h	fef44703	;
assign	mem[11'd1051]	=	32'h	00d00793	;
assign	mem[11'd1052]	=	32'h	00f71a63	;
assign	mem[11'd1053]	=	32'h	00000517	;
assign	mem[11'd1054]	=	32'h	06850513	;
assign	mem[11'd1055]	=	32'h	f51ff0ef	;
assign	mem[11'd1056]	=	32'h	0100006f	;
assign	mem[11'd1057]	=	32'h	fef44783	;
assign	mem[11'd1058]	=	32'h	00078513	;
assign	mem[11'd1059]	=	32'h	ef9ff0ef	;
assign	mem[11'd1060]	=	32'h	fef44783	;
assign	mem[11'd1061]	=	32'h	00078513	;
assign	mem[11'd1062]	=	32'h	01c12083	;
assign	mem[11'd1063]	=	32'h	01812403	;
assign	mem[11'd1064]	=	32'h	02010113	;
assign	mem[11'd1065]	=	32'h	00008067	;
assign	mem[11'd1066]	=	32'h	00000a0d	;
assign	mem[11'd1067]	=	32'h	20636f73	;
assign	mem[11'd1068]	=	32'h	0000203e	;
assign	mem[11'd1069]	=	32'h	00000d20	;
assign	mem[11'd1070]	=	32'h	656c6966	;
assign	mem[11'd1071]	=	32'h	00000000	;
assign	mem[11'd1072]	=	32'h	0000006a	;
assign	mem[11'd1073]	=	32'h	00000070	;
assign	mem[11'd1074]	=	32'h	00000069	;
assign	mem[11'd1075]	=	32'h	6e550d0a	;
assign	mem[11'd1076]	=	32'h	776f6e6b	;
assign	mem[11'd1077]	=	32'h	00203a6e	;
assign	mem[11'd1078]	=	32'h	00000d0a	;
assign	mem[11'd1079]	=	32'h	00000a0d	;
           
endmodule

module bios_mem_test (
    input clk,
    input ena,
    input rst,
    input [10:0] addra,
    output reg [31:0] douta,
    input enb,
    input [10:0] addrb,
    output reg [31:0] doutb
);

    wire [31:0] mem [2048-1:0];
    always @(posedge clk) begin
        if (rst) begin
            douta <= 32'b0;
        end
        else if (ena) begin
            douta <= mem[addra];
        end
    end

    always @(posedge clk) begin
        if (rst) begin
            doutb <= 32'b0;
        end
        else if (enb) begin
            doutb <= mem[addrb];
        end
    end
//machine code for demo bios
    assign mem[11'd0000] = 32'h00000013;
    assign mem[11'd0001] = 32'h00000013;
    assign mem[11'd0002] = 32'h00000013;
    assign mem[11'd0003] = 32'h00000013;
    assign mem[11'd0004] = 32'h00000013;
    assign mem[11'd0005] = 32'h10000fb7;
    assign mem[11'd0006] = 32'h000f8067;
    assign mem[11'd0007] = 32'h00000013;
    assign mem[11'd0008] = 32'h00000013;
    assign mem[11'd0009] = 32'h00000013;
    assign mem[11'd0010] = 32'h00000013;
    assign mem[11'd0011] = 32'h00000013;

endmodule