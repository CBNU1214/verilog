`timescale 1 ps / 1 ps

(* RESET_PC = "1073741824" *) 
(* STRUCTURAL_NETLIST = "yes" *)
module RISCV_TOP_netlist
   (CLK,
    RSTn,
    I_MEM_CSN,
    I_MEM_DOUT,
    I_MEM_ADDR,
    D_MEM_CSN,
    D_MEM_DOUT,
    D_MEM_DI,
    D_MEM_ADDR,
    D_MEM_WEN,
    D_MEM_BE,
    RF_WE,
    RF_RA1,
    RF_RA2,
    RF_WA,
    RF_RD1,
    RF_RD2,
    RF_WD,
    CRF_WE,
    CRF_RA1,
    CRF_RA2,
    CRF_WA,
    CRF_RD1,
    CRF_RD2,
    CRF_WD);
  input CLK;
  input RSTn;
  output I_MEM_CSN;
  input [31:0]I_MEM_DOUT;
  output [31:0]I_MEM_ADDR;
  output D_MEM_CSN;
  input [31:0]D_MEM_DOUT;
  output [31:0]D_MEM_DI;
  output [31:0]D_MEM_ADDR;
  output D_MEM_WEN;
  output [3:0]D_MEM_BE;
  output RF_WE;
  output [4:0]RF_RA1;
  output [4:0]RF_RA2;
  output [4:0]RF_WA;
  input [31:0]RF_RD1;
  input [31:0]RF_RD2;
  output [31:0]RF_WD;
  output CRF_WE;
  output [4:0]CRF_RA1;
  output [4:0]CRF_RA2;
  output [4:0]CRF_WA;
  input [31:0]CRF_RD1;
  input [31:0]CRF_RD2;
  output [31:0]CRF_WD;

  wire \<const0> ;
  wire \<const1> ;
  wire [31:0]ALU_DIN1;
  wire [31:0]ALU_DIN2;
  wire CLK;
  wire CLK_IBUF;
  wire CLK_IBUF_BUFG;
  wire [4:0]CRF_RA1;
  wire [4:0]CRF_RA1_OBUF;
  wire [4:0]CRF_RA2;
  wire [4:0]CRF_RA2_OBUF;
  wire [31:0]CRF_RD1;
  wire [31:0]CRF_RD1_IBUF;
  wire [31:0]CRF_RD2;
  wire [31:0]CRF_RD2_IBUF;
  wire [4:0]CRF_WA;
  wire [4:0]CRF_WA_OBUF;
  wire [31:0]CRF_WD;
  wire [31:0]CRF_WD_OBUF;
  wire CRF_WE;
  wire CRF_WE_OBUF;
  wire [31:0]CUSTOM_ALU_OUT;
  wire [31:26]CUSTOM_ALU_SEL;
  wire CUSTOM_EN;
  wire [2:1]CUSTOM_INSTRUCTION_STALL_CYCLE;
  wire CUSTOM_RD;
  wire CUSTOM_RS1;
  wire CUSTOM_RS2;
  wire [30:30]D0;
  wire [29:0]DECODED_INSTRUCTION;
  wire [2:0]DIN1_FORWARD;
  wire [2:0]DIN2_FORWARD;
  wire [31:0]D_MEM_ADDR;
  wire [31:0]D_MEM_ADDR_OBUF;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_13_n_1 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_13_n_2 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_13_n_3 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_15_n_1 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_15_n_2 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_15_n_3 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_21_n_1 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_21_n_2 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_21_n_3 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_24_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_25_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_26_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_26_n_1 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_26_n_2 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_26_n_3 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_27_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_28_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_29_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_30_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_31_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_32_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_33_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_34_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[0]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[10]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_9_n_1 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_9_n_2 ;
  wire \D_MEM_ADDR_OBUF[11]_inst_i_9_n_3 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[12]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[13]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[14]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_24_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_25_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_26_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_27_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_28_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_29_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_30_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_31_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_32_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_33_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[15]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[16]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[17]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[18]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[19]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[1]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[20]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[21]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[22]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_24_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_25_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_26_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_27_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_28_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_29_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[23]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[24]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[25]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[27]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_6_n_1 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_6_n_2 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_6_n_3 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[28]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[29]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[2]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[30]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_24_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_25_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_26_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_27_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_28_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_29_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_30_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_31_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_32_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_33_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_34_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_35_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_5_n_2 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_5_n_3 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_6_n_1 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_6_n_2 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_6_n_3 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_7_n_1 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_7_n_2 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_7_n_3 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[31]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_24_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_25_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_26_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_27_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_28_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_29_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_30_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_31_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_32_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_9_n_1 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_9_n_2 ;
  wire \D_MEM_ADDR_OBUF[3]_inst_i_9_n_3 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[4]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[5]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[6]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_22_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_23_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_24_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_25_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_26_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_27_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_9_n_1 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_9_n_2 ;
  wire \D_MEM_ADDR_OBUF[7]_inst_i_9_n_3 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_8_n_1 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_8_n_2 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_8_n_3 ;
  wire \D_MEM_ADDR_OBUF[8]_inst_i_9_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_10_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_11_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_12_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_13_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_14_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_15_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_16_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_17_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_18_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_19_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_20_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_21_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_2_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_3_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_4_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_5_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_6_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_7_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_8_n_0 ;
  wire \D_MEM_ADDR_OBUF[9]_inst_i_9_n_0 ;
  wire [3:0]D_MEM_BE;
  wire [3:0]D_MEM_BE_OBUF;
  wire D_MEM_CSN;
  wire D_MEM_CSN_OBUF;
  wire [31:0]D_MEM_DI;
  wire [31:0]D_MEM_DI_OBUF;
  wire [31:0]D_MEM_DOUT;
  wire [31:0]D_MEM_DOUT_IBUF;
  wire D_MEM_WEN;
  wire D_MEM_WEN_OBUF;
  wire EX_BR_TAKEN;
  wire [31:26]EX_CUSTOM_ALU_SEL;
  wire EX_CUSTOM_RD;
  wire [39:0]EX_MEM_Q;
  wire [31:0]EX_RF_RD1;
  wire [31:0]EX_RF_RD2;
  wire \FF_CUSTOM_EN/Q_reg_n_0_[0] ;
  wire \FF_EX_MEM_TEMP/Q_reg_n_0_[0] ;
  wire \FF_EX_MEM_TEMP/Q_reg_n_0_[1] ;
  wire \FF_ID_EX/Q_reg[158]_rep__0_n_0 ;
  wire \FF_ID_EX/Q_reg[158]_rep__1_n_0 ;
  wire \FF_ID_EX/Q_reg[158]_rep__2_n_0 ;
  wire \FF_ID_EX/Q_reg[158]_rep__3_n_0 ;
  wire \FF_ID_EX/Q_reg[158]_rep__4_n_0 ;
  wire \FF_ID_EX/Q_reg[158]_rep_n_0 ;
  wire \FF_ID_EX/Q_reg[170]_rep__0_n_0 ;
  wire \FF_ID_EX/Q_reg[170]_rep__1_n_0 ;
  wire \FF_ID_EX/Q_reg[170]_rep__2_n_0 ;
  wire \FF_ID_EX/Q_reg[170]_rep__3_n_0 ;
  wire \FF_ID_EX/Q_reg[170]_rep_n_0 ;
  wire \FF_ID_EX/Q_reg_n_0_[158] ;
  wire \FF_ID_EX/Q_reg_n_0_[164] ;
  wire \FF_ID_EX/Q_reg_n_0_[165] ;
  wire \FF_ID_EX/Q_reg_n_0_[168] ;
  wire \FF_ID_EX/Q_reg_n_0_[169] ;
  wire \FF_ID_EX/Q_reg_n_0_[170] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[0] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[10] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[11] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[12] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[13] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[14] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[15] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[16] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[17] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[18] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[19] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[1] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[20] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[21] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[22] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[23] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[24] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[25] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[26] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[27] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[28] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[29] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[2] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[30] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[31] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[3] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[4] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[5] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[6] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[7] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[8] ;
  wire \FF_IF_ID_PCADD/Q_reg_n_0_[9] ;
  wire \FF_JALR_EN/Q_reg_n_0_[0] ;
  wire GND_2;
  wire ID_BR;
  wire [171:112]ID_EX_D;
  wire [161:0]ID_EX_Q;
  wire [31:0]ID_IMMEDIATE;
  wire ID_IMMEDIATE_EN;
  wire ID_JAL_AFTER_LU;
  wire ID_MEM;
  wire [31:0]ID_PC;
  wire [31:0]ID_RD2_FORWARDED;
  wire ID_WB_AFTER_LU;
  wire ID_WE_AFTER_LU3;
  wire [31:0]IF_PC2;
  wire [31:1]IF_PC_ADD4;
  wire INT0_carry__0_i_10_n_0;
  wire INT0_carry__0_i_11_n_0;
  wire INT0_carry__0_i_12_n_0;
  wire INT0_carry__0_i_13_n_0;
  wire INT0_carry__0_i_14_n_0;
  wire INT0_carry__0_i_15_n_0;
  wire INT0_carry__0_i_16_n_0;
  wire INT0_carry__0_i_17_n_0;
  wire INT0_carry__0_i_18_n_0;
  wire INT0_carry__0_i_19_n_0;
  wire INT0_carry__0_i_20_n_0;
  wire INT0_carry__0_i_21_n_0;
  wire INT0_carry__0_i_22_n_0;
  wire INT0_carry__0_i_23_n_0;
  wire INT0_carry__0_i_5_n_0;
  wire INT0_carry__0_i_6_n_0;
  wire INT0_carry__0_i_7_n_0;
  wire INT0_carry__0_i_8_n_0;
  wire INT0_carry__0_i_9_n_0;
  wire INT0_carry__1_i_10_n_0;
  wire INT0_carry__1_i_11_n_0;
  wire INT0_carry__1_i_12_n_0;
  wire INT0_carry__1_i_13_n_0;
  wire INT0_carry__1_i_14_n_0;
  wire INT0_carry__1_i_2_n_0;
  wire INT0_carry__1_i_5_n_0;
  wire INT0_carry__1_i_6_n_0;
  wire INT0_carry__1_i_7_n_0;
  wire INT0_carry__1_i_8_n_0;
  wire INT0_carry__1_i_9_n_0;
  wire INT0_carry__2_i_10_n_0;
  wire INT0_carry__2_i_11_n_0;
  wire INT0_carry__2_i_12_n_0;
  wire INT0_carry__2_i_13_n_0;
  wire INT0_carry__2_i_14_n_0;
  wire INT0_carry__2_i_15_n_0;
  wire INT0_carry__2_i_16_n_0;
  wire INT0_carry__2_i_1_n_0;
  wire INT0_carry__2_i_2_n_0;
  wire INT0_carry__2_i_5_n_0;
  wire INT0_carry__2_i_6_n_0;
  wire INT0_carry__2_i_7_n_0;
  wire INT0_carry__2_i_8_n_0;
  wire INT0_carry__2_i_9_n_0;
  wire INT0_carry__3_i_1_n_0;
  wire INT0_carry__3_i_2_n_0;
  wire INT0_carry__3_i_3_n_0;
  wire INT0_carry__3_i_4_n_0;
  wire INT0_carry__3_i_5_n_0;
  wire INT0_carry__3_i_6_n_0;
  wire INT0_carry__3_i_7_n_0;
  wire INT0_carry__3_i_8_n_0;
  wire INT0_carry__4_i_2_n_0;
  wire INT0_carry__4_i_4_n_0;
  wire INT0_carry__4_i_5_n_0;
  wire INT0_carry__4_i_6_n_0;
  wire INT0_carry_i_10_n_0;
  wire INT0_carry_i_11_n_0;
  wire INT0_carry_i_12_n_0;
  wire INT0_carry_i_13_n_0;
  wire INT0_carry_i_14_n_0;
  wire INT0_carry_i_15_n_0;
  wire INT0_carry_i_16_n_0;
  wire INT0_carry_i_17_n_0;
  wire INT0_carry_i_18_n_0;
  wire INT0_carry_i_19_n_0;
  wire INT0_carry_i_20_n_0;
  wire INT0_carry_i_21_n_0;
  wire INT0_carry_i_22_n_0;
  wire INT0_carry_i_23_n_0;
  wire INT0_carry_i_24_n_0;
  wire INT0_carry_i_25_n_0;
  wire INT0_carry_i_26_n_0;
  wire INT0_carry_i_27_n_0;
  wire INT0_carry_i_28_n_0;
  wire INT0_carry_i_29_n_0;
  wire INT0_carry_i_6_n_0;
  wire INT0_carry_i_7_n_0;
  wire INT0_carry_i_8_n_0;
  wire INT0_carry_i_9_n_0;
  wire [31:0]I_MEM_ADDR;
  wire [31:0]I_MEM_ADDR_OBUF;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_2_n_0 ;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_2_n_1 ;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_2_n_2 ;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_2_n_3 ;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_3_n_0 ;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_4_n_0 ;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[11]_inst_i_6_n_0 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_2_n_0 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_2_n_1 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_2_n_2 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_2_n_3 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_3_n_0 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_4_n_0 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[15]_inst_i_6_n_0 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_2_n_0 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_2_n_1 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_2_n_2 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_2_n_3 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_3_n_0 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_4_n_0 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[19]_inst_i_6_n_0 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_2_n_0 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_2_n_1 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_2_n_2 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_2_n_3 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_3_n_0 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_4_n_0 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[23]_inst_i_6_n_0 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_2_n_0 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_2_n_1 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_2_n_2 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_2_n_3 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_3_n_0 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_4_n_0 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[27]_inst_i_6_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_10_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_12_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_3_n_1 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_3_n_2 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_3_n_3 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_4_n_1 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_4_n_2 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_4_n_3 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_6_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_7_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_8_n_0 ;
  wire \I_MEM_ADDR_OBUF[31]_inst_i_9_n_0 ;
  wire \I_MEM_ADDR_OBUF[3]_inst_i_2_n_0 ;
  wire \I_MEM_ADDR_OBUF[3]_inst_i_2_n_1 ;
  wire \I_MEM_ADDR_OBUF[3]_inst_i_2_n_2 ;
  wire \I_MEM_ADDR_OBUF[3]_inst_i_2_n_3 ;
  wire \I_MEM_ADDR_OBUF[3]_inst_i_3_n_0 ;
  wire \I_MEM_ADDR_OBUF[3]_inst_i_4_n_0 ;
  wire \I_MEM_ADDR_OBUF[3]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_2_n_0 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_2_n_1 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_2_n_2 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_2_n_3 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_3_n_0 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_4_n_0 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_5_n_0 ;
  wire \I_MEM_ADDR_OBUF[7]_inst_i_6_n_0 ;
  wire I_MEM_CSN;
  wire [31:0]I_MEM_DOUT;
  wire [11:2]I_MEM_DOUT_FILTERED;
  wire [31:2]I_MEM_DOUT_IBUF;
  wire LU_HAZARD;
  wire MEM_CUSTOM_RD;
  wire MEM_D_MEM_ALU_FINAL1;
  wire [6:1]MEM_LOAD_SEL;
  wire [37:37]MEM_WB_Q;
  wire PSUM0__0_carry__0_i_10__0_n_0;
  wire PSUM0__0_carry__0_i_10__1_n_0;
  wire PSUM0__0_carry__0_i_10__2_n_0;
  wire PSUM0__0_carry__0_i_10_n_0;
  wire PSUM0__0_carry__0_i_11__0_n_0;
  wire PSUM0__0_carry__0_i_11__1_n_0;
  wire PSUM0__0_carry__0_i_11__2_n_0;
  wire PSUM0__0_carry__0_i_11_n_0;
  wire PSUM0__0_carry__0_i_12__0_n_0;
  wire PSUM0__0_carry__0_i_12__1_n_0;
  wire PSUM0__0_carry__0_i_12__2_n_0;
  wire PSUM0__0_carry__0_i_12_n_0;
  wire PSUM0__0_carry__0_i_1__0_n_0;
  wire PSUM0__0_carry__0_i_1__1_n_0;
  wire PSUM0__0_carry__0_i_1__2_n_0;
  wire PSUM0__0_carry__0_i_1_n_0;
  wire PSUM0__0_carry__0_i_2__0_n_0;
  wire PSUM0__0_carry__0_i_2__1_n_0;
  wire PSUM0__0_carry__0_i_2__2_n_0;
  wire PSUM0__0_carry__0_i_2_n_0;
  wire PSUM0__0_carry__0_i_3__0_n_0;
  wire PSUM0__0_carry__0_i_3__1_n_0;
  wire PSUM0__0_carry__0_i_3__2_n_0;
  wire PSUM0__0_carry__0_i_3_n_0;
  wire PSUM0__0_carry__0_i_4__0_n_0;
  wire PSUM0__0_carry__0_i_4__1_n_0;
  wire PSUM0__0_carry__0_i_4__2_n_0;
  wire PSUM0__0_carry__0_i_4_n_0;
  wire PSUM0__0_carry__0_i_5__0_n_0;
  wire PSUM0__0_carry__0_i_5__1_n_0;
  wire PSUM0__0_carry__0_i_5__2_n_0;
  wire PSUM0__0_carry__0_i_5_n_0;
  wire PSUM0__0_carry__0_i_6__0_n_0;
  wire PSUM0__0_carry__0_i_6__1_n_0;
  wire PSUM0__0_carry__0_i_6__2_n_0;
  wire PSUM0__0_carry__0_i_6_n_0;
  wire PSUM0__0_carry__0_i_7__0_n_0;
  wire PSUM0__0_carry__0_i_7__1_n_0;
  wire PSUM0__0_carry__0_i_7__2_n_0;
  wire PSUM0__0_carry__0_i_7_n_0;
  wire PSUM0__0_carry__0_i_8__0_n_0;
  wire PSUM0__0_carry__0_i_8__1_n_0;
  wire PSUM0__0_carry__0_i_8__2_n_0;
  wire PSUM0__0_carry__0_i_8_n_0;
  wire PSUM0__0_carry__0_i_9__0_n_0;
  wire PSUM0__0_carry__0_i_9__1_n_0;
  wire PSUM0__0_carry__0_i_9__2_n_0;
  wire PSUM0__0_carry__0_i_9_n_0;
  wire PSUM0__0_carry__1_i_1__0_n_0;
  wire PSUM0__0_carry__1_i_1__1_n_0;
  wire PSUM0__0_carry__1_i_1__2_n_0;
  wire PSUM0__0_carry__1_i_1_n_0;
  wire PSUM0__0_carry__1_i_2__0_n_0;
  wire PSUM0__0_carry__1_i_2__1_n_0;
  wire PSUM0__0_carry__1_i_2__2_n_0;
  wire PSUM0__0_carry__1_i_2_n_0;
  wire PSUM0__0_carry__1_i_3__0_n_0;
  wire PSUM0__0_carry__1_i_3__1_n_0;
  wire PSUM0__0_carry__1_i_3__2_n_0;
  wire PSUM0__0_carry__1_i_3_n_0;
  wire PSUM0__0_carry__1_i_4__0_n_0;
  wire PSUM0__0_carry__1_i_4__1_n_0;
  wire PSUM0__0_carry__1_i_4__2_n_0;
  wire PSUM0__0_carry__1_i_4_n_0;
  wire PSUM0__0_carry_i_1__0_n_0;
  wire PSUM0__0_carry_i_1__1_n_0;
  wire PSUM0__0_carry_i_1__2_n_0;
  wire PSUM0__0_carry_i_1_n_0;
  wire PSUM0__0_carry_i_2__0_n_0;
  wire PSUM0__0_carry_i_2__1_n_0;
  wire PSUM0__0_carry_i_2__2_n_0;
  wire PSUM0__0_carry_i_2_n_0;
  wire PSUM0__0_carry_i_3__0_n_0;
  wire PSUM0__0_carry_i_3__1_n_0;
  wire PSUM0__0_carry_i_3__2_n_0;
  wire PSUM0__0_carry_i_3_n_0;
  wire PSUM0__0_carry_i_4__0_n_0;
  wire PSUM0__0_carry_i_4__1_n_0;
  wire PSUM0__0_carry_i_4__2_n_0;
  wire PSUM0__0_carry_i_4_n_0;
  wire PSUM0__0_carry_i_5__0_n_0;
  wire PSUM0__0_carry_i_5__1_n_0;
  wire PSUM0__0_carry_i_5__2_n_0;
  wire PSUM0__0_carry_i_5_n_0;
  wire PSUM0__0_carry_i_6__0_n_0;
  wire PSUM0__0_carry_i_6__1_n_0;
  wire PSUM0__0_carry_i_6__2_n_0;
  wire PSUM0__0_carry_i_6_n_0;
  wire PSUM0__0_carry_i_7__0_n_0;
  wire PSUM0__0_carry_i_7__1_n_0;
  wire PSUM0__0_carry_i_7__2_n_0;
  wire PSUM0__0_carry_i_7_n_0;
  wire PSUM0__0_carry_i_8__0_n_0;
  wire PSUM0__0_carry_i_8__1_n_0;
  wire PSUM0__0_carry_i_8__2_n_0;
  wire PSUM0__0_carry_i_8_n_0;
  wire PSUM0__30_carry__0_i_10__0_n_0;
  wire PSUM0__30_carry__0_i_10__1_n_0;
  wire PSUM0__30_carry__0_i_10__2_n_0;
  wire PSUM0__30_carry__0_i_10_n_0;
  wire PSUM0__30_carry__0_i_11__0_n_0;
  wire PSUM0__30_carry__0_i_11__1_n_0;
  wire PSUM0__30_carry__0_i_11__2_n_0;
  wire PSUM0__30_carry__0_i_11_n_0;
  wire PSUM0__30_carry__0_i_12__0_n_0;
  wire PSUM0__30_carry__0_i_12__1_n_0;
  wire PSUM0__30_carry__0_i_12__2_n_0;
  wire PSUM0__30_carry__0_i_12_n_0;
  wire PSUM0__30_carry__0_i_1__0_n_0;
  wire PSUM0__30_carry__0_i_1__1_n_0;
  wire PSUM0__30_carry__0_i_1__2_n_0;
  wire PSUM0__30_carry__0_i_1_n_0;
  wire PSUM0__30_carry__0_i_2__0_n_0;
  wire PSUM0__30_carry__0_i_2__1_n_0;
  wire PSUM0__30_carry__0_i_2__2_n_0;
  wire PSUM0__30_carry__0_i_2_n_0;
  wire PSUM0__30_carry__0_i_3__0_n_0;
  wire PSUM0__30_carry__0_i_3__1_n_0;
  wire PSUM0__30_carry__0_i_3__2_n_0;
  wire PSUM0__30_carry__0_i_3_n_0;
  wire PSUM0__30_carry__0_i_4__0_n_0;
  wire PSUM0__30_carry__0_i_4__1_n_0;
  wire PSUM0__30_carry__0_i_4__2_n_0;
  wire PSUM0__30_carry__0_i_4_n_0;
  wire PSUM0__30_carry__0_i_5__0_n_0;
  wire PSUM0__30_carry__0_i_5__1_n_0;
  wire PSUM0__30_carry__0_i_5__2_n_0;
  wire PSUM0__30_carry__0_i_5_n_0;
  wire PSUM0__30_carry__0_i_6__0_n_0;
  wire PSUM0__30_carry__0_i_6__1_n_0;
  wire PSUM0__30_carry__0_i_6__2_n_0;
  wire PSUM0__30_carry__0_i_6_n_0;
  wire PSUM0__30_carry__0_i_7__0_n_0;
  wire PSUM0__30_carry__0_i_7__1_n_0;
  wire PSUM0__30_carry__0_i_7__2_n_0;
  wire PSUM0__30_carry__0_i_7_n_0;
  wire PSUM0__30_carry__0_i_8__0_n_0;
  wire PSUM0__30_carry__0_i_8__1_n_0;
  wire PSUM0__30_carry__0_i_8__2_n_0;
  wire PSUM0__30_carry__0_i_8_n_0;
  wire PSUM0__30_carry__0_i_9__0_n_0;
  wire PSUM0__30_carry__0_i_9__1_n_0;
  wire PSUM0__30_carry__0_i_9__2_n_0;
  wire PSUM0__30_carry__0_i_9_n_0;
  wire PSUM0__30_carry__1_i_1__0_n_0;
  wire PSUM0__30_carry__1_i_1__1_n_0;
  wire PSUM0__30_carry__1_i_1__2_n_0;
  wire PSUM0__30_carry__1_i_1_n_0;
  wire PSUM0__30_carry__1_i_2__0_n_0;
  wire PSUM0__30_carry__1_i_2__1_n_0;
  wire PSUM0__30_carry__1_i_2__2_n_0;
  wire PSUM0__30_carry__1_i_2_n_0;
  wire PSUM0__30_carry__1_i_3__0_n_0;
  wire PSUM0__30_carry__1_i_3__1_n_0;
  wire PSUM0__30_carry__1_i_3__2_n_0;
  wire PSUM0__30_carry__1_i_3_n_0;
  wire PSUM0__30_carry__1_i_4__0_n_0;
  wire PSUM0__30_carry__1_i_4__1_n_0;
  wire PSUM0__30_carry__1_i_4__2_n_0;
  wire PSUM0__30_carry__1_i_4_n_0;
  wire PSUM0__30_carry_i_1__0_n_0;
  wire PSUM0__30_carry_i_1__1_n_0;
  wire PSUM0__30_carry_i_1__2_n_0;
  wire PSUM0__30_carry_i_1_n_0;
  wire PSUM0__30_carry_i_2__0_n_0;
  wire PSUM0__30_carry_i_2__1_n_0;
  wire PSUM0__30_carry_i_2__2_n_0;
  wire PSUM0__30_carry_i_2_n_0;
  wire PSUM0__30_carry_i_3__0_n_0;
  wire PSUM0__30_carry_i_3__1_n_0;
  wire PSUM0__30_carry_i_3__2_n_0;
  wire PSUM0__30_carry_i_3_n_0;
  wire PSUM0__30_carry_i_4__0_n_0;
  wire PSUM0__30_carry_i_4__1_n_0;
  wire PSUM0__30_carry_i_4__2_n_0;
  wire PSUM0__30_carry_i_4_n_0;
  wire PSUM0__30_carry_i_5__0_n_0;
  wire PSUM0__30_carry_i_5__1_n_0;
  wire PSUM0__30_carry_i_5__2_n_0;
  wire PSUM0__30_carry_i_5_n_0;
  wire PSUM0__30_carry_i_6__0_n_0;
  wire PSUM0__30_carry_i_6__1_n_0;
  wire PSUM0__30_carry_i_6__2_n_0;
  wire PSUM0__30_carry_i_6_n_0;
  wire PSUM0__30_carry_i_7__0_n_0;
  wire PSUM0__30_carry_i_7__1_n_0;
  wire PSUM0__30_carry_i_7__2_n_0;
  wire PSUM0__30_carry_i_7_n_0;
  wire PSUM0__30_carry_i_8__0_n_0;
  wire PSUM0__30_carry_i_8__1_n_0;
  wire PSUM0__30_carry_i_8__2_n_0;
  wire PSUM0__30_carry_i_8_n_0;
  wire PSUM0__60_carry__0_i_10__0_n_0;
  wire PSUM0__60_carry__0_i_10__1_n_0;
  wire PSUM0__60_carry__0_i_10__2_n_0;
  wire PSUM0__60_carry__0_i_10_n_0;
  wire PSUM0__60_carry__0_i_11__0_n_0;
  wire PSUM0__60_carry__0_i_11__1_n_0;
  wire PSUM0__60_carry__0_i_11__2_n_0;
  wire PSUM0__60_carry__0_i_11_n_0;
  wire PSUM0__60_carry__0_i_12__0_n_0;
  wire PSUM0__60_carry__0_i_12__1_n_0;
  wire PSUM0__60_carry__0_i_12__2_n_0;
  wire PSUM0__60_carry__0_i_12_n_0;
  wire PSUM0__60_carry__0_i_13__0_n_0;
  wire PSUM0__60_carry__0_i_13__1_n_0;
  wire PSUM0__60_carry__0_i_13__2_n_0;
  wire PSUM0__60_carry__0_i_13_n_0;
  wire PSUM0__60_carry__0_i_14__0_n_0;
  wire PSUM0__60_carry__0_i_14__1_n_0;
  wire PSUM0__60_carry__0_i_14__2_n_0;
  wire PSUM0__60_carry__0_i_14_n_0;
  wire PSUM0__60_carry__0_i_15__0_n_0;
  wire PSUM0__60_carry__0_i_15__1_n_0;
  wire PSUM0__60_carry__0_i_15__2_n_0;
  wire PSUM0__60_carry__0_i_15_n_0;
  wire PSUM0__60_carry__0_i_1__0_n_0;
  wire PSUM0__60_carry__0_i_1__1_n_0;
  wire PSUM0__60_carry__0_i_1__2_n_0;
  wire PSUM0__60_carry__0_i_1_n_0;
  wire PSUM0__60_carry__0_i_2__0_n_0;
  wire PSUM0__60_carry__0_i_2__1_n_0;
  wire PSUM0__60_carry__0_i_2__2_n_0;
  wire PSUM0__60_carry__0_i_2_n_0;
  wire PSUM0__60_carry__0_i_3__0_n_0;
  wire PSUM0__60_carry__0_i_3__1_n_0;
  wire PSUM0__60_carry__0_i_3__2_n_0;
  wire PSUM0__60_carry__0_i_3_n_0;
  wire PSUM0__60_carry__0_i_4__0_n_0;
  wire PSUM0__60_carry__0_i_4__1_n_0;
  wire PSUM0__60_carry__0_i_4__2_n_0;
  wire PSUM0__60_carry__0_i_4_n_0;
  wire PSUM0__60_carry__0_i_5__0_n_0;
  wire PSUM0__60_carry__0_i_5__1_n_0;
  wire PSUM0__60_carry__0_i_5__2_n_0;
  wire PSUM0__60_carry__0_i_5_n_0;
  wire PSUM0__60_carry__0_i_6__0_n_0;
  wire PSUM0__60_carry__0_i_6__1_n_0;
  wire PSUM0__60_carry__0_i_6__2_n_0;
  wire PSUM0__60_carry__0_i_6_n_0;
  wire PSUM0__60_carry__0_i_7__0_n_0;
  wire PSUM0__60_carry__0_i_7__1_n_0;
  wire PSUM0__60_carry__0_i_7__2_n_0;
  wire PSUM0__60_carry__0_i_7_n_0;
  wire PSUM0__60_carry__0_i_8__0_n_0;
  wire PSUM0__60_carry__0_i_8__1_n_0;
  wire PSUM0__60_carry__0_i_8__2_n_0;
  wire PSUM0__60_carry__0_i_8_n_0;
  wire PSUM0__60_carry__0_i_9__0_n_0;
  wire PSUM0__60_carry__0_i_9__1_n_0;
  wire PSUM0__60_carry__0_i_9__2_n_0;
  wire PSUM0__60_carry__0_i_9_n_0;
  wire PSUM0__60_carry__1_i_10__0_n_0;
  wire PSUM0__60_carry__1_i_10__1_n_0;
  wire PSUM0__60_carry__1_i_10__2_n_0;
  wire PSUM0__60_carry__1_i_10_n_0;
  wire PSUM0__60_carry__1_i_11__0_n_0;
  wire PSUM0__60_carry__1_i_11__1_n_0;
  wire PSUM0__60_carry__1_i_11__2_n_0;
  wire PSUM0__60_carry__1_i_11_n_0;
  wire PSUM0__60_carry__1_i_12__0_n_0;
  wire PSUM0__60_carry__1_i_12__1_n_0;
  wire PSUM0__60_carry__1_i_12__2_n_0;
  wire PSUM0__60_carry__1_i_12_n_0;
  wire PSUM0__60_carry__1_i_13__0_n_0;
  wire PSUM0__60_carry__1_i_13__1_n_0;
  wire PSUM0__60_carry__1_i_13__2_n_0;
  wire PSUM0__60_carry__1_i_13_n_0;
  wire PSUM0__60_carry__1_i_14__0_n_0;
  wire PSUM0__60_carry__1_i_14__1_n_0;
  wire PSUM0__60_carry__1_i_14__2_n_0;
  wire PSUM0__60_carry__1_i_14_n_0;
  wire PSUM0__60_carry__1_i_15__0_n_0;
  wire PSUM0__60_carry__1_i_15__1_n_0;
  wire PSUM0__60_carry__1_i_15__2_n_0;
  wire PSUM0__60_carry__1_i_15_n_0;
  wire PSUM0__60_carry__1_i_1__0_n_0;
  wire PSUM0__60_carry__1_i_1__1_n_0;
  wire PSUM0__60_carry__1_i_1__2_n_0;
  wire PSUM0__60_carry__1_i_1_n_0;
  wire PSUM0__60_carry__1_i_2__0_n_0;
  wire PSUM0__60_carry__1_i_2__1_n_0;
  wire PSUM0__60_carry__1_i_2__2_n_0;
  wire PSUM0__60_carry__1_i_2_n_0;
  wire PSUM0__60_carry__1_i_3__0_n_0;
  wire PSUM0__60_carry__1_i_3__1_n_0;
  wire PSUM0__60_carry__1_i_3__2_n_0;
  wire PSUM0__60_carry__1_i_3_n_0;
  wire PSUM0__60_carry__1_i_4__0_n_0;
  wire PSUM0__60_carry__1_i_4__1_n_0;
  wire PSUM0__60_carry__1_i_4__2_n_0;
  wire PSUM0__60_carry__1_i_4_n_0;
  wire PSUM0__60_carry__1_i_5__0_n_0;
  wire PSUM0__60_carry__1_i_5__1_n_0;
  wire PSUM0__60_carry__1_i_5__2_n_0;
  wire PSUM0__60_carry__1_i_5_n_0;
  wire PSUM0__60_carry__1_i_6__0_n_0;
  wire PSUM0__60_carry__1_i_6__1_n_0;
  wire PSUM0__60_carry__1_i_6__2_n_0;
  wire PSUM0__60_carry__1_i_6_n_0;
  wire PSUM0__60_carry__1_i_7__0_n_0;
  wire PSUM0__60_carry__1_i_7__1_n_0;
  wire PSUM0__60_carry__1_i_7__2_n_0;
  wire PSUM0__60_carry__1_i_7_n_0;
  wire PSUM0__60_carry__1_i_8__0_n_0;
  wire PSUM0__60_carry__1_i_8__1_n_0;
  wire PSUM0__60_carry__1_i_8__2_n_0;
  wire PSUM0__60_carry__1_i_8_n_0;
  wire PSUM0__60_carry__1_i_9__0_n_0;
  wire PSUM0__60_carry__1_i_9__1_n_0;
  wire PSUM0__60_carry__1_i_9__2_n_0;
  wire PSUM0__60_carry__1_i_9_n_0;
  wire PSUM0__60_carry__2_i_1__0_n_0;
  wire PSUM0__60_carry__2_i_1__1_n_0;
  wire PSUM0__60_carry__2_i_1__2_n_0;
  wire PSUM0__60_carry__2_i_1_n_0;
  wire PSUM0__60_carry_i_1__0_n_0;
  wire PSUM0__60_carry_i_1__1_n_0;
  wire PSUM0__60_carry_i_1__2_n_0;
  wire PSUM0__60_carry_i_1_n_0;
  wire PSUM0__60_carry_i_2__0_n_0;
  wire PSUM0__60_carry_i_2__1_n_0;
  wire PSUM0__60_carry_i_2__2_n_0;
  wire PSUM0__60_carry_i_2_n_0;
  wire PSUM0__60_carry_i_3__0_n_0;
  wire PSUM0__60_carry_i_3__1_n_0;
  wire PSUM0__60_carry_i_3__2_n_0;
  wire PSUM0__60_carry_i_3_n_0;
  wire PSUM0__60_carry_i_4__0_n_0;
  wire PSUM0__60_carry_i_4__1_n_0;
  wire PSUM0__60_carry_i_4__2_n_0;
  wire PSUM0__60_carry_i_4_n_0;
  wire PSUM0__60_carry_i_5__0_n_0;
  wire PSUM0__60_carry_i_5__1_n_0;
  wire PSUM0__60_carry_i_5__2_n_0;
  wire PSUM0__60_carry_i_5_n_0;
  wire PSUM1__0_carry__0_i_10__0_n_0;
  wire PSUM1__0_carry__0_i_10__1_n_0;
  wire PSUM1__0_carry__0_i_10_n_0;
  wire PSUM1__0_carry__0_i_11__0_n_0;
  wire PSUM1__0_carry__0_i_11__1_n_0;
  wire PSUM1__0_carry__0_i_11__2_n_0;
  wire PSUM1__0_carry__0_i_11_n_0;
  wire PSUM1__0_carry__0_i_12__0_n_0;
  wire PSUM1__0_carry__0_i_12__1_n_0;
  wire PSUM1__0_carry__0_i_12__2_n_0;
  wire PSUM1__0_carry__0_i_12_n_0;
  wire PSUM1__0_carry__0_i_13_n_0;
  wire PSUM1__0_carry__0_i_1__0_n_0;
  wire PSUM1__0_carry__0_i_1__1_n_0;
  wire PSUM1__0_carry__0_i_1__2_n_0;
  wire PSUM1__0_carry__0_i_1_n_0;
  wire PSUM1__0_carry__0_i_2__0_n_0;
  wire PSUM1__0_carry__0_i_2__1_n_0;
  wire PSUM1__0_carry__0_i_2__2_n_0;
  wire PSUM1__0_carry__0_i_2_n_0;
  wire PSUM1__0_carry__0_i_3__0_n_0;
  wire PSUM1__0_carry__0_i_3__1_n_0;
  wire PSUM1__0_carry__0_i_3__2_n_0;
  wire PSUM1__0_carry__0_i_3_n_0;
  wire PSUM1__0_carry__0_i_4__0_n_0;
  wire PSUM1__0_carry__0_i_4__1_n_0;
  wire PSUM1__0_carry__0_i_4__2_n_0;
  wire PSUM1__0_carry__0_i_4_n_0;
  wire PSUM1__0_carry__0_i_5__0_n_0;
  wire PSUM1__0_carry__0_i_5__1_n_0;
  wire PSUM1__0_carry__0_i_5__2_n_0;
  wire PSUM1__0_carry__0_i_5_n_0;
  wire PSUM1__0_carry__0_i_6__0_n_0;
  wire PSUM1__0_carry__0_i_6__1_n_0;
  wire PSUM1__0_carry__0_i_6__2_n_0;
  wire PSUM1__0_carry__0_i_6_n_0;
  wire PSUM1__0_carry__0_i_7__0_n_0;
  wire PSUM1__0_carry__0_i_7__1_n_0;
  wire PSUM1__0_carry__0_i_7__2_n_0;
  wire PSUM1__0_carry__0_i_7_n_0;
  wire PSUM1__0_carry__0_i_8__0_n_0;
  wire PSUM1__0_carry__0_i_8__1_n_0;
  wire PSUM1__0_carry__0_i_8__2_n_0;
  wire PSUM1__0_carry__0_i_8_n_0;
  wire PSUM1__0_carry__0_i_9__0_n_0;
  wire PSUM1__0_carry__0_i_9__1_n_0;
  wire PSUM1__0_carry__0_i_9__2_n_0;
  wire PSUM1__0_carry__0_i_9_n_0;
  wire PSUM1__0_carry__1_i_1__0_n_0;
  wire PSUM1__0_carry__1_i_1__1_n_0;
  wire PSUM1__0_carry__1_i_1__2_n_0;
  wire PSUM1__0_carry__1_i_1_n_0;
  wire PSUM1__0_carry__1_i_2__0_n_0;
  wire PSUM1__0_carry__1_i_2__1_n_0;
  wire PSUM1__0_carry__1_i_2__2_n_0;
  wire PSUM1__0_carry__1_i_2_n_0;
  wire PSUM1__0_carry__1_i_3__0_n_0;
  wire PSUM1__0_carry__1_i_3__1_n_0;
  wire PSUM1__0_carry__1_i_3__2_n_0;
  wire PSUM1__0_carry__1_i_3_n_0;
  wire PSUM1__0_carry__1_i_4__0_n_0;
  wire PSUM1__0_carry__1_i_4__1_n_0;
  wire PSUM1__0_carry__1_i_4__2_n_0;
  wire PSUM1__0_carry__1_i_4_n_0;
  wire PSUM1__0_carry_i_1__0_n_0;
  wire PSUM1__0_carry_i_1__1_n_0;
  wire PSUM1__0_carry_i_1__2_n_0;
  wire PSUM1__0_carry_i_1_n_0;
  wire PSUM1__0_carry_i_2__0_n_0;
  wire PSUM1__0_carry_i_2__1_n_0;
  wire PSUM1__0_carry_i_2__2_n_0;
  wire PSUM1__0_carry_i_2_n_0;
  wire PSUM1__0_carry_i_3__0_n_0;
  wire PSUM1__0_carry_i_3__1_n_0;
  wire PSUM1__0_carry_i_3__2_n_0;
  wire PSUM1__0_carry_i_3_n_0;
  wire PSUM1__0_carry_i_4__0_n_0;
  wire PSUM1__0_carry_i_4__1_n_0;
  wire PSUM1__0_carry_i_4__2_n_0;
  wire PSUM1__0_carry_i_4_n_0;
  wire PSUM1__0_carry_i_5__0_n_0;
  wire PSUM1__0_carry_i_5__1_n_0;
  wire PSUM1__0_carry_i_5__2_n_0;
  wire PSUM1__0_carry_i_5_n_0;
  wire PSUM1__0_carry_i_6__0_n_0;
  wire PSUM1__0_carry_i_6__1_n_0;
  wire PSUM1__0_carry_i_6__2_n_0;
  wire PSUM1__0_carry_i_6_n_0;
  wire PSUM1__0_carry_i_7__0_n_0;
  wire PSUM1__0_carry_i_7__1_n_0;
  wire PSUM1__0_carry_i_7__2_n_0;
  wire PSUM1__0_carry_i_7_n_0;
  wire PSUM1__0_carry_i_8__0_n_0;
  wire PSUM1__0_carry_i_8__1_n_0;
  wire PSUM1__0_carry_i_8__2_n_0;
  wire PSUM1__0_carry_i_8_n_0;
  wire PSUM1__30_carry__0_i_10__0_n_0;
  wire PSUM1__30_carry__0_i_10__1_n_0;
  wire PSUM1__30_carry__0_i_10__2_n_0;
  wire PSUM1__30_carry__0_i_10_n_0;
  wire PSUM1__30_carry__0_i_11__0_n_0;
  wire PSUM1__30_carry__0_i_11__1_n_0;
  wire PSUM1__30_carry__0_i_11__2_n_0;
  wire PSUM1__30_carry__0_i_11_n_0;
  wire PSUM1__30_carry__0_i_12__0_n_0;
  wire PSUM1__30_carry__0_i_12__1_n_0;
  wire PSUM1__30_carry__0_i_12__2_n_0;
  wire PSUM1__30_carry__0_i_12_n_0;
  wire PSUM1__30_carry__0_i_1__0_n_0;
  wire PSUM1__30_carry__0_i_1__1_n_0;
  wire PSUM1__30_carry__0_i_1__2_n_0;
  wire PSUM1__30_carry__0_i_1_n_0;
  wire PSUM1__30_carry__0_i_2__0_n_0;
  wire PSUM1__30_carry__0_i_2__1_n_0;
  wire PSUM1__30_carry__0_i_2__2_n_0;
  wire PSUM1__30_carry__0_i_2_n_0;
  wire PSUM1__30_carry__0_i_3__0_n_0;
  wire PSUM1__30_carry__0_i_3__1_n_0;
  wire PSUM1__30_carry__0_i_3__2_n_0;
  wire PSUM1__30_carry__0_i_3_n_0;
  wire PSUM1__30_carry__0_i_4__0_n_0;
  wire PSUM1__30_carry__0_i_4__1_n_0;
  wire PSUM1__30_carry__0_i_4__2_n_0;
  wire PSUM1__30_carry__0_i_4_n_0;
  wire PSUM1__30_carry__0_i_5__0_n_0;
  wire PSUM1__30_carry__0_i_5__1_n_0;
  wire PSUM1__30_carry__0_i_5__2_n_0;
  wire PSUM1__30_carry__0_i_5_n_0;
  wire PSUM1__30_carry__0_i_6__0_n_0;
  wire PSUM1__30_carry__0_i_6__1_n_0;
  wire PSUM1__30_carry__0_i_6__2_n_0;
  wire PSUM1__30_carry__0_i_6_n_0;
  wire PSUM1__30_carry__0_i_7__0_n_0;
  wire PSUM1__30_carry__0_i_7__1_n_0;
  wire PSUM1__30_carry__0_i_7__2_n_0;
  wire PSUM1__30_carry__0_i_7_n_0;
  wire PSUM1__30_carry__0_i_8__0_n_0;
  wire PSUM1__30_carry__0_i_8__1_n_0;
  wire PSUM1__30_carry__0_i_8__2_n_0;
  wire PSUM1__30_carry__0_i_8_n_0;
  wire PSUM1__30_carry__0_i_9__0_n_0;
  wire PSUM1__30_carry__0_i_9__1_n_0;
  wire PSUM1__30_carry__0_i_9__2_n_0;
  wire PSUM1__30_carry__0_i_9_n_0;
  wire PSUM1__30_carry__1_i_1__0_n_0;
  wire PSUM1__30_carry__1_i_1__1_n_0;
  wire PSUM1__30_carry__1_i_1__2_n_0;
  wire PSUM1__30_carry__1_i_1_n_0;
  wire PSUM1__30_carry__1_i_2__0_n_0;
  wire PSUM1__30_carry__1_i_2__1_n_0;
  wire PSUM1__30_carry__1_i_2__2_n_0;
  wire PSUM1__30_carry__1_i_2_n_0;
  wire PSUM1__30_carry__1_i_3__0_n_0;
  wire PSUM1__30_carry__1_i_3__1_n_0;
  wire PSUM1__30_carry__1_i_3__2_n_0;
  wire PSUM1__30_carry__1_i_3_n_0;
  wire PSUM1__30_carry__1_i_4__0_n_0;
  wire PSUM1__30_carry__1_i_4__1_n_0;
  wire PSUM1__30_carry__1_i_4__2_n_0;
  wire PSUM1__30_carry__1_i_4_n_0;
  wire PSUM1__30_carry_i_1__0_n_0;
  wire PSUM1__30_carry_i_1__1_n_0;
  wire PSUM1__30_carry_i_1__2_n_0;
  wire PSUM1__30_carry_i_1_n_0;
  wire PSUM1__30_carry_i_2__0_n_0;
  wire PSUM1__30_carry_i_2__1_n_0;
  wire PSUM1__30_carry_i_2__2_n_0;
  wire PSUM1__30_carry_i_2_n_0;
  wire PSUM1__30_carry_i_3__0_n_0;
  wire PSUM1__30_carry_i_3__1_n_0;
  wire PSUM1__30_carry_i_3__2_n_0;
  wire PSUM1__30_carry_i_3_n_0;
  wire PSUM1__30_carry_i_4__0_n_0;
  wire PSUM1__30_carry_i_4__1_n_0;
  wire PSUM1__30_carry_i_4__2_n_0;
  wire PSUM1__30_carry_i_4_n_0;
  wire PSUM1__30_carry_i_5__0_n_0;
  wire PSUM1__30_carry_i_5__1_n_0;
  wire PSUM1__30_carry_i_5__2_n_0;
  wire PSUM1__30_carry_i_5_n_0;
  wire PSUM1__30_carry_i_6__0_n_0;
  wire PSUM1__30_carry_i_6__1_n_0;
  wire PSUM1__30_carry_i_6__2_n_0;
  wire PSUM1__30_carry_i_6_n_0;
  wire PSUM1__30_carry_i_7__0_n_0;
  wire PSUM1__30_carry_i_7__1_n_0;
  wire PSUM1__30_carry_i_7__2_n_0;
  wire PSUM1__30_carry_i_7_n_0;
  wire PSUM1__30_carry_i_8__0_n_0;
  wire PSUM1__30_carry_i_8__1_n_0;
  wire PSUM1__30_carry_i_8__2_n_0;
  wire PSUM1__30_carry_i_8_n_0;
  wire PSUM1__60_carry__0_i_10__0_n_0;
  wire PSUM1__60_carry__0_i_10__1_n_0;
  wire PSUM1__60_carry__0_i_10__2_n_0;
  wire PSUM1__60_carry__0_i_10_n_0;
  wire PSUM1__60_carry__0_i_11__0_n_0;
  wire PSUM1__60_carry__0_i_11__1_n_0;
  wire PSUM1__60_carry__0_i_11__2_n_0;
  wire PSUM1__60_carry__0_i_11_n_0;
  wire PSUM1__60_carry__0_i_12__0_n_0;
  wire PSUM1__60_carry__0_i_12__1_n_0;
  wire PSUM1__60_carry__0_i_12__2_n_0;
  wire PSUM1__60_carry__0_i_12_n_0;
  wire PSUM1__60_carry__0_i_13__0_n_0;
  wire PSUM1__60_carry__0_i_13__1_n_0;
  wire PSUM1__60_carry__0_i_13__2_n_0;
  wire PSUM1__60_carry__0_i_13_n_0;
  wire PSUM1__60_carry__0_i_14__0_n_0;
  wire PSUM1__60_carry__0_i_14__1_n_0;
  wire PSUM1__60_carry__0_i_14__2_n_0;
  wire PSUM1__60_carry__0_i_14_n_0;
  wire PSUM1__60_carry__0_i_15__0_n_0;
  wire PSUM1__60_carry__0_i_15__1_n_0;
  wire PSUM1__60_carry__0_i_15__2_n_0;
  wire PSUM1__60_carry__0_i_15_n_0;
  wire PSUM1__60_carry__0_i_1__0_n_0;
  wire PSUM1__60_carry__0_i_1__1_n_0;
  wire PSUM1__60_carry__0_i_1__2_n_0;
  wire PSUM1__60_carry__0_i_1_n_0;
  wire PSUM1__60_carry__0_i_2__0_n_0;
  wire PSUM1__60_carry__0_i_2__1_n_0;
  wire PSUM1__60_carry__0_i_2__2_n_0;
  wire PSUM1__60_carry__0_i_2_n_0;
  wire PSUM1__60_carry__0_i_3__0_n_0;
  wire PSUM1__60_carry__0_i_3__1_n_0;
  wire PSUM1__60_carry__0_i_3__2_n_0;
  wire PSUM1__60_carry__0_i_3_n_0;
  wire PSUM1__60_carry__0_i_4__0_n_0;
  wire PSUM1__60_carry__0_i_4__1_n_0;
  wire PSUM1__60_carry__0_i_4__2_n_0;
  wire PSUM1__60_carry__0_i_4_n_0;
  wire PSUM1__60_carry__0_i_5__0_n_0;
  wire PSUM1__60_carry__0_i_5__1_n_0;
  wire PSUM1__60_carry__0_i_5__2_n_0;
  wire PSUM1__60_carry__0_i_5_n_0;
  wire PSUM1__60_carry__0_i_6__0_n_0;
  wire PSUM1__60_carry__0_i_6__1_n_0;
  wire PSUM1__60_carry__0_i_6__2_n_0;
  wire PSUM1__60_carry__0_i_6_n_0;
  wire PSUM1__60_carry__0_i_7__0_n_0;
  wire PSUM1__60_carry__0_i_7__1_n_0;
  wire PSUM1__60_carry__0_i_7__2_n_0;
  wire PSUM1__60_carry__0_i_7_n_0;
  wire PSUM1__60_carry__0_i_8__0_n_0;
  wire PSUM1__60_carry__0_i_8__1_n_0;
  wire PSUM1__60_carry__0_i_8__2_n_0;
  wire PSUM1__60_carry__0_i_8_n_0;
  wire PSUM1__60_carry__0_i_9__0_n_0;
  wire PSUM1__60_carry__0_i_9__1_n_0;
  wire PSUM1__60_carry__0_i_9__2_n_0;
  wire PSUM1__60_carry__0_i_9_n_0;
  wire PSUM1__60_carry__1_i_10__0_n_0;
  wire PSUM1__60_carry__1_i_10__1_n_0;
  wire PSUM1__60_carry__1_i_10__2_n_0;
  wire PSUM1__60_carry__1_i_10_n_0;
  wire PSUM1__60_carry__1_i_11__0_n_0;
  wire PSUM1__60_carry__1_i_11__1_n_0;
  wire PSUM1__60_carry__1_i_11__2_n_0;
  wire PSUM1__60_carry__1_i_11_n_0;
  wire PSUM1__60_carry__1_i_12__0_n_0;
  wire PSUM1__60_carry__1_i_12__1_n_0;
  wire PSUM1__60_carry__1_i_12__2_n_0;
  wire PSUM1__60_carry__1_i_12_n_0;
  wire PSUM1__60_carry__1_i_13__0_n_0;
  wire PSUM1__60_carry__1_i_13__1_n_0;
  wire PSUM1__60_carry__1_i_13__2_n_0;
  wire PSUM1__60_carry__1_i_13_n_0;
  wire PSUM1__60_carry__1_i_14__0_n_0;
  wire PSUM1__60_carry__1_i_14__1_n_0;
  wire PSUM1__60_carry__1_i_14__2_n_0;
  wire PSUM1__60_carry__1_i_14_n_0;
  wire PSUM1__60_carry__1_i_15__0_n_0;
  wire PSUM1__60_carry__1_i_15__1_n_0;
  wire PSUM1__60_carry__1_i_15__2_n_0;
  wire PSUM1__60_carry__1_i_15_n_0;
  wire PSUM1__60_carry__1_i_1__0_n_0;
  wire PSUM1__60_carry__1_i_1__1_n_0;
  wire PSUM1__60_carry__1_i_1__2_n_0;
  wire PSUM1__60_carry__1_i_1_n_0;
  wire PSUM1__60_carry__1_i_2__0_n_0;
  wire PSUM1__60_carry__1_i_2__1_n_0;
  wire PSUM1__60_carry__1_i_2__2_n_0;
  wire PSUM1__60_carry__1_i_2_n_0;
  wire PSUM1__60_carry__1_i_3__0_n_0;
  wire PSUM1__60_carry__1_i_3__1_n_0;
  wire PSUM1__60_carry__1_i_3__2_n_0;
  wire PSUM1__60_carry__1_i_3_n_0;
  wire PSUM1__60_carry__1_i_4__0_n_0;
  wire PSUM1__60_carry__1_i_4__1_n_0;
  wire PSUM1__60_carry__1_i_4__2_n_0;
  wire PSUM1__60_carry__1_i_4_n_0;
  wire PSUM1__60_carry__1_i_5__0_n_0;
  wire PSUM1__60_carry__1_i_5__1_n_0;
  wire PSUM1__60_carry__1_i_5__2_n_0;
  wire PSUM1__60_carry__1_i_5_n_0;
  wire PSUM1__60_carry__1_i_6__0_n_0;
  wire PSUM1__60_carry__1_i_6__1_n_0;
  wire PSUM1__60_carry__1_i_6__2_n_0;
  wire PSUM1__60_carry__1_i_6_n_0;
  wire PSUM1__60_carry__1_i_7__0_n_0;
  wire PSUM1__60_carry__1_i_7__1_n_0;
  wire PSUM1__60_carry__1_i_7__2_n_0;
  wire PSUM1__60_carry__1_i_7_n_0;
  wire PSUM1__60_carry__1_i_8__0_n_0;
  wire PSUM1__60_carry__1_i_8__1_n_0;
  wire PSUM1__60_carry__1_i_8__2_n_0;
  wire PSUM1__60_carry__1_i_8_n_0;
  wire PSUM1__60_carry__1_i_9__0_n_0;
  wire PSUM1__60_carry__1_i_9__1_n_0;
  wire PSUM1__60_carry__1_i_9__2_n_0;
  wire PSUM1__60_carry__1_i_9_n_0;
  wire PSUM1__60_carry__2_i_1__0_n_0;
  wire PSUM1__60_carry__2_i_1__1_n_0;
  wire PSUM1__60_carry__2_i_1__2_n_0;
  wire PSUM1__60_carry__2_i_1_n_0;
  wire PSUM1__60_carry_i_1__0_n_0;
  wire PSUM1__60_carry_i_1__1_n_0;
  wire PSUM1__60_carry_i_1__2_n_0;
  wire PSUM1__60_carry_i_1_n_0;
  wire PSUM1__60_carry_i_2__0_n_0;
  wire PSUM1__60_carry_i_2__1_n_0;
  wire PSUM1__60_carry_i_2__2_n_0;
  wire PSUM1__60_carry_i_2_n_0;
  wire PSUM1__60_carry_i_3__0_n_0;
  wire PSUM1__60_carry_i_3__1_n_0;
  wire PSUM1__60_carry_i_3__2_n_0;
  wire PSUM1__60_carry_i_3_n_0;
  wire PSUM1__60_carry_i_4__0_n_0;
  wire PSUM1__60_carry_i_4__1_n_0;
  wire PSUM1__60_carry_i_4__2_n_0;
  wire PSUM1__60_carry_i_4_n_0;
  wire PSUM1__60_carry_i_5__0_n_0;
  wire PSUM1__60_carry_i_5__1_n_0;
  wire PSUM1__60_carry_i_5__2_n_0;
  wire PSUM1__60_carry_i_5_n_0;
  wire PSUM2__0_carry__0_i_10__0_n_0;
  wire PSUM2__0_carry__0_i_10__1_n_0;
  wire PSUM2__0_carry__0_i_10__2_n_0;
  wire PSUM2__0_carry__0_i_10_n_0;
  wire PSUM2__0_carry__0_i_11__0_n_0;
  wire PSUM2__0_carry__0_i_11__1_n_0;
  wire PSUM2__0_carry__0_i_11__2_n_0;
  wire PSUM2__0_carry__0_i_11_n_0;
  wire PSUM2__0_carry__0_i_12__0_n_0;
  wire PSUM2__0_carry__0_i_12__1_n_0;
  wire PSUM2__0_carry__0_i_12__2_n_0;
  wire PSUM2__0_carry__0_i_12_n_0;
  wire PSUM2__0_carry__0_i_1__0_n_0;
  wire PSUM2__0_carry__0_i_1__1_n_0;
  wire PSUM2__0_carry__0_i_1__2_n_0;
  wire PSUM2__0_carry__0_i_1_n_0;
  wire PSUM2__0_carry__0_i_2__0_n_0;
  wire PSUM2__0_carry__0_i_2__1_n_0;
  wire PSUM2__0_carry__0_i_2__2_n_0;
  wire PSUM2__0_carry__0_i_2_n_0;
  wire PSUM2__0_carry__0_i_3__0_n_0;
  wire PSUM2__0_carry__0_i_3__1_n_0;
  wire PSUM2__0_carry__0_i_3__2_n_0;
  wire PSUM2__0_carry__0_i_3_n_0;
  wire PSUM2__0_carry__0_i_4__0_n_0;
  wire PSUM2__0_carry__0_i_4__1_n_0;
  wire PSUM2__0_carry__0_i_4__2_n_0;
  wire PSUM2__0_carry__0_i_4_n_0;
  wire PSUM2__0_carry__0_i_5__0_n_0;
  wire PSUM2__0_carry__0_i_5__1_n_0;
  wire PSUM2__0_carry__0_i_5__2_n_0;
  wire PSUM2__0_carry__0_i_5_n_0;
  wire PSUM2__0_carry__0_i_6__0_n_0;
  wire PSUM2__0_carry__0_i_6__1_n_0;
  wire PSUM2__0_carry__0_i_6__2_n_0;
  wire PSUM2__0_carry__0_i_6_n_0;
  wire PSUM2__0_carry__0_i_7__0_n_0;
  wire PSUM2__0_carry__0_i_7__1_n_0;
  wire PSUM2__0_carry__0_i_7__2_n_0;
  wire PSUM2__0_carry__0_i_7_n_0;
  wire PSUM2__0_carry__0_i_8__0_n_0;
  wire PSUM2__0_carry__0_i_8__1_n_0;
  wire PSUM2__0_carry__0_i_8__2_n_0;
  wire PSUM2__0_carry__0_i_8_n_0;
  wire PSUM2__0_carry__0_i_9__0_n_0;
  wire PSUM2__0_carry__0_i_9__1_n_0;
  wire PSUM2__0_carry__0_i_9__2_n_0;
  wire PSUM2__0_carry__0_i_9_n_0;
  wire PSUM2__0_carry__1_i_1__0_n_0;
  wire PSUM2__0_carry__1_i_1__1_n_0;
  wire PSUM2__0_carry__1_i_1__2_n_0;
  wire PSUM2__0_carry__1_i_1_n_0;
  wire PSUM2__0_carry__1_i_2__0_n_0;
  wire PSUM2__0_carry__1_i_2__1_n_0;
  wire PSUM2__0_carry__1_i_2__2_n_0;
  wire PSUM2__0_carry__1_i_2_n_0;
  wire PSUM2__0_carry__1_i_3__0_n_0;
  wire PSUM2__0_carry__1_i_3__1_n_0;
  wire PSUM2__0_carry__1_i_3__2_n_0;
  wire PSUM2__0_carry__1_i_3_n_0;
  wire PSUM2__0_carry__1_i_4__0_n_0;
  wire PSUM2__0_carry__1_i_4__1_n_0;
  wire PSUM2__0_carry__1_i_4__2_n_0;
  wire PSUM2__0_carry__1_i_4_n_0;
  wire PSUM2__0_carry_i_1__0_n_0;
  wire PSUM2__0_carry_i_1__1_n_0;
  wire PSUM2__0_carry_i_1__2_n_0;
  wire PSUM2__0_carry_i_1_n_0;
  wire PSUM2__0_carry_i_2__0_n_0;
  wire PSUM2__0_carry_i_2__1_n_0;
  wire PSUM2__0_carry_i_2__2_n_0;
  wire PSUM2__0_carry_i_2_n_0;
  wire PSUM2__0_carry_i_3__0_n_0;
  wire PSUM2__0_carry_i_3__1_n_0;
  wire PSUM2__0_carry_i_3__2_n_0;
  wire PSUM2__0_carry_i_3_n_0;
  wire PSUM2__0_carry_i_4__0_n_0;
  wire PSUM2__0_carry_i_4__1_n_0;
  wire PSUM2__0_carry_i_4__2_n_0;
  wire PSUM2__0_carry_i_4_n_0;
  wire PSUM2__0_carry_i_5__0_n_0;
  wire PSUM2__0_carry_i_5__1_n_0;
  wire PSUM2__0_carry_i_5__2_n_0;
  wire PSUM2__0_carry_i_5_n_0;
  wire PSUM2__0_carry_i_6__0_n_0;
  wire PSUM2__0_carry_i_6__1_n_0;
  wire PSUM2__0_carry_i_6__2_n_0;
  wire PSUM2__0_carry_i_6_n_0;
  wire PSUM2__0_carry_i_7__0_n_0;
  wire PSUM2__0_carry_i_7__1_n_0;
  wire PSUM2__0_carry_i_7__2_n_0;
  wire PSUM2__0_carry_i_7_n_0;
  wire PSUM2__0_carry_i_8__0_n_0;
  wire PSUM2__0_carry_i_8__1_n_0;
  wire PSUM2__0_carry_i_8__2_n_0;
  wire PSUM2__0_carry_i_8_n_0;
  wire PSUM2__30_carry__0_i_10__0_n_0;
  wire PSUM2__30_carry__0_i_10__1_n_0;
  wire PSUM2__30_carry__0_i_10__2_n_0;
  wire PSUM2__30_carry__0_i_10_n_0;
  wire PSUM2__30_carry__0_i_11__0_n_0;
  wire PSUM2__30_carry__0_i_11__1_n_0;
  wire PSUM2__30_carry__0_i_11__2_n_0;
  wire PSUM2__30_carry__0_i_11_n_0;
  wire PSUM2__30_carry__0_i_12__0_n_0;
  wire PSUM2__30_carry__0_i_12__1_n_0;
  wire PSUM2__30_carry__0_i_12__2_n_0;
  wire PSUM2__30_carry__0_i_12_n_0;
  wire PSUM2__30_carry__0_i_1__0_n_0;
  wire PSUM2__30_carry__0_i_1__1_n_0;
  wire PSUM2__30_carry__0_i_1__2_n_0;
  wire PSUM2__30_carry__0_i_1_n_0;
  wire PSUM2__30_carry__0_i_2__0_n_0;
  wire PSUM2__30_carry__0_i_2__1_n_0;
  wire PSUM2__30_carry__0_i_2__2_n_0;
  wire PSUM2__30_carry__0_i_2_n_0;
  wire PSUM2__30_carry__0_i_3__0_n_0;
  wire PSUM2__30_carry__0_i_3__1_n_0;
  wire PSUM2__30_carry__0_i_3__2_n_0;
  wire PSUM2__30_carry__0_i_3_n_0;
  wire PSUM2__30_carry__0_i_4__0_n_0;
  wire PSUM2__30_carry__0_i_4__1_n_0;
  wire PSUM2__30_carry__0_i_4__2_n_0;
  wire PSUM2__30_carry__0_i_4_n_0;
  wire PSUM2__30_carry__0_i_5__0_n_0;
  wire PSUM2__30_carry__0_i_5__1_n_0;
  wire PSUM2__30_carry__0_i_5__2_n_0;
  wire PSUM2__30_carry__0_i_5_n_0;
  wire PSUM2__30_carry__0_i_6__0_n_0;
  wire PSUM2__30_carry__0_i_6__1_n_0;
  wire PSUM2__30_carry__0_i_6__2_n_0;
  wire PSUM2__30_carry__0_i_6_n_0;
  wire PSUM2__30_carry__0_i_7__0_n_0;
  wire PSUM2__30_carry__0_i_7__1_n_0;
  wire PSUM2__30_carry__0_i_7__2_n_0;
  wire PSUM2__30_carry__0_i_7_n_0;
  wire PSUM2__30_carry__0_i_8__0_n_0;
  wire PSUM2__30_carry__0_i_8__1_n_0;
  wire PSUM2__30_carry__0_i_8__2_n_0;
  wire PSUM2__30_carry__0_i_8_n_0;
  wire PSUM2__30_carry__0_i_9__0_n_0;
  wire PSUM2__30_carry__0_i_9__1_n_0;
  wire PSUM2__30_carry__0_i_9__2_n_0;
  wire PSUM2__30_carry__0_i_9_n_0;
  wire PSUM2__30_carry__1_i_1__0_n_0;
  wire PSUM2__30_carry__1_i_1__1_n_0;
  wire PSUM2__30_carry__1_i_1__2_n_0;
  wire PSUM2__30_carry__1_i_1_n_0;
  wire PSUM2__30_carry__1_i_2__0_n_0;
  wire PSUM2__30_carry__1_i_2__1_n_0;
  wire PSUM2__30_carry__1_i_2__2_n_0;
  wire PSUM2__30_carry__1_i_2_n_0;
  wire PSUM2__30_carry__1_i_3__0_n_0;
  wire PSUM2__30_carry__1_i_3__1_n_0;
  wire PSUM2__30_carry__1_i_3__2_n_0;
  wire PSUM2__30_carry__1_i_3_n_0;
  wire PSUM2__30_carry__1_i_4__0_n_0;
  wire PSUM2__30_carry__1_i_4__1_n_0;
  wire PSUM2__30_carry__1_i_4__2_n_0;
  wire PSUM2__30_carry__1_i_4_n_0;
  wire PSUM2__30_carry_i_1__0_n_0;
  wire PSUM2__30_carry_i_1__1_n_0;
  wire PSUM2__30_carry_i_1__2_n_0;
  wire PSUM2__30_carry_i_1_n_0;
  wire PSUM2__30_carry_i_2__0_n_0;
  wire PSUM2__30_carry_i_2__1_n_0;
  wire PSUM2__30_carry_i_2__2_n_0;
  wire PSUM2__30_carry_i_2_n_0;
  wire PSUM2__30_carry_i_3__0_n_0;
  wire PSUM2__30_carry_i_3__1_n_0;
  wire PSUM2__30_carry_i_3__2_n_0;
  wire PSUM2__30_carry_i_3_n_0;
  wire PSUM2__30_carry_i_4__0_n_0;
  wire PSUM2__30_carry_i_4__1_n_0;
  wire PSUM2__30_carry_i_4__2_n_0;
  wire PSUM2__30_carry_i_4_n_0;
  wire PSUM2__30_carry_i_5__0_n_0;
  wire PSUM2__30_carry_i_5__1_n_0;
  wire PSUM2__30_carry_i_5__2_n_0;
  wire PSUM2__30_carry_i_5_n_0;
  wire PSUM2__30_carry_i_6__0_n_0;
  wire PSUM2__30_carry_i_6__1_n_0;
  wire PSUM2__30_carry_i_6__2_n_0;
  wire PSUM2__30_carry_i_6_n_0;
  wire PSUM2__30_carry_i_7__0_n_0;
  wire PSUM2__30_carry_i_7__1_n_0;
  wire PSUM2__30_carry_i_7__2_n_0;
  wire PSUM2__30_carry_i_7_n_0;
  wire PSUM2__30_carry_i_8__0_n_0;
  wire PSUM2__30_carry_i_8__1_n_0;
  wire PSUM2__30_carry_i_8__2_n_0;
  wire PSUM2__30_carry_i_8_n_0;
  wire PSUM2__60_carry__0_i_10__0_n_0;
  wire PSUM2__60_carry__0_i_10__1_n_0;
  wire PSUM2__60_carry__0_i_10__2_n_0;
  wire PSUM2__60_carry__0_i_10_n_0;
  wire PSUM2__60_carry__0_i_11__0_n_0;
  wire PSUM2__60_carry__0_i_11__1_n_0;
  wire PSUM2__60_carry__0_i_11__2_n_0;
  wire PSUM2__60_carry__0_i_11_n_0;
  wire PSUM2__60_carry__0_i_12__0_n_0;
  wire PSUM2__60_carry__0_i_12__1_n_0;
  wire PSUM2__60_carry__0_i_12__2_n_0;
  wire PSUM2__60_carry__0_i_12_n_0;
  wire PSUM2__60_carry__0_i_13__0_n_0;
  wire PSUM2__60_carry__0_i_13__1_n_0;
  wire PSUM2__60_carry__0_i_13__2_n_0;
  wire PSUM2__60_carry__0_i_13_n_0;
  wire PSUM2__60_carry__0_i_14__0_n_0;
  wire PSUM2__60_carry__0_i_14__1_n_0;
  wire PSUM2__60_carry__0_i_14__2_n_0;
  wire PSUM2__60_carry__0_i_14_n_0;
  wire PSUM2__60_carry__0_i_15__0_n_0;
  wire PSUM2__60_carry__0_i_15__1_n_0;
  wire PSUM2__60_carry__0_i_15__2_n_0;
  wire PSUM2__60_carry__0_i_15_n_0;
  wire PSUM2__60_carry__0_i_1__0_n_0;
  wire PSUM2__60_carry__0_i_1__1_n_0;
  wire PSUM2__60_carry__0_i_1__2_n_0;
  wire PSUM2__60_carry__0_i_1_n_0;
  wire PSUM2__60_carry__0_i_2__0_n_0;
  wire PSUM2__60_carry__0_i_2__1_n_0;
  wire PSUM2__60_carry__0_i_2__2_n_0;
  wire PSUM2__60_carry__0_i_2_n_0;
  wire PSUM2__60_carry__0_i_3__0_n_0;
  wire PSUM2__60_carry__0_i_3__1_n_0;
  wire PSUM2__60_carry__0_i_3__2_n_0;
  wire PSUM2__60_carry__0_i_3_n_0;
  wire PSUM2__60_carry__0_i_4__0_n_0;
  wire PSUM2__60_carry__0_i_4__1_n_0;
  wire PSUM2__60_carry__0_i_4__2_n_0;
  wire PSUM2__60_carry__0_i_4_n_0;
  wire PSUM2__60_carry__0_i_5__0_n_0;
  wire PSUM2__60_carry__0_i_5__1_n_0;
  wire PSUM2__60_carry__0_i_5__2_n_0;
  wire PSUM2__60_carry__0_i_5_n_0;
  wire PSUM2__60_carry__0_i_6__0_n_0;
  wire PSUM2__60_carry__0_i_6__1_n_0;
  wire PSUM2__60_carry__0_i_6__2_n_0;
  wire PSUM2__60_carry__0_i_6_n_0;
  wire PSUM2__60_carry__0_i_7__0_n_0;
  wire PSUM2__60_carry__0_i_7__1_n_0;
  wire PSUM2__60_carry__0_i_7__2_n_0;
  wire PSUM2__60_carry__0_i_7_n_0;
  wire PSUM2__60_carry__0_i_8__0_n_0;
  wire PSUM2__60_carry__0_i_8__1_n_0;
  wire PSUM2__60_carry__0_i_8__2_n_0;
  wire PSUM2__60_carry__0_i_8_n_0;
  wire PSUM2__60_carry__0_i_9__0_n_0;
  wire PSUM2__60_carry__0_i_9__1_n_0;
  wire PSUM2__60_carry__0_i_9__2_n_0;
  wire PSUM2__60_carry__0_i_9_n_0;
  wire PSUM2__60_carry__1_i_10__0_n_0;
  wire PSUM2__60_carry__1_i_10__1_n_0;
  wire PSUM2__60_carry__1_i_10__2_n_0;
  wire PSUM2__60_carry__1_i_10_n_0;
  wire PSUM2__60_carry__1_i_11__0_n_0;
  wire PSUM2__60_carry__1_i_11__1_n_0;
  wire PSUM2__60_carry__1_i_11__2_n_0;
  wire PSUM2__60_carry__1_i_11_n_0;
  wire PSUM2__60_carry__1_i_12__0_n_0;
  wire PSUM2__60_carry__1_i_12__1_n_0;
  wire PSUM2__60_carry__1_i_12__2_n_0;
  wire PSUM2__60_carry__1_i_12_n_0;
  wire PSUM2__60_carry__1_i_13__0_n_0;
  wire PSUM2__60_carry__1_i_13__1_n_0;
  wire PSUM2__60_carry__1_i_13__2_n_0;
  wire PSUM2__60_carry__1_i_13_n_0;
  wire PSUM2__60_carry__1_i_14__0_n_0;
  wire PSUM2__60_carry__1_i_14__1_n_0;
  wire PSUM2__60_carry__1_i_14__2_n_0;
  wire PSUM2__60_carry__1_i_14_n_0;
  wire PSUM2__60_carry__1_i_15__0_n_0;
  wire PSUM2__60_carry__1_i_15__1_n_0;
  wire PSUM2__60_carry__1_i_15__2_n_0;
  wire PSUM2__60_carry__1_i_15_n_0;
  wire PSUM2__60_carry__1_i_1__0_n_0;
  wire PSUM2__60_carry__1_i_1__1_n_0;
  wire PSUM2__60_carry__1_i_1__2_n_0;
  wire PSUM2__60_carry__1_i_1_n_0;
  wire PSUM2__60_carry__1_i_2__0_n_0;
  wire PSUM2__60_carry__1_i_2__1_n_0;
  wire PSUM2__60_carry__1_i_2__2_n_0;
  wire PSUM2__60_carry__1_i_2_n_0;
  wire PSUM2__60_carry__1_i_3__0_n_0;
  wire PSUM2__60_carry__1_i_3__1_n_0;
  wire PSUM2__60_carry__1_i_3__2_n_0;
  wire PSUM2__60_carry__1_i_3_n_0;
  wire PSUM2__60_carry__1_i_4__0_n_0;
  wire PSUM2__60_carry__1_i_4__1_n_0;
  wire PSUM2__60_carry__1_i_4__2_n_0;
  wire PSUM2__60_carry__1_i_4_n_0;
  wire PSUM2__60_carry__1_i_5__0_n_0;
  wire PSUM2__60_carry__1_i_5__1_n_0;
  wire PSUM2__60_carry__1_i_5__2_n_0;
  wire PSUM2__60_carry__1_i_5_n_0;
  wire PSUM2__60_carry__1_i_6__0_n_0;
  wire PSUM2__60_carry__1_i_6__1_n_0;
  wire PSUM2__60_carry__1_i_6__2_n_0;
  wire PSUM2__60_carry__1_i_6_n_0;
  wire PSUM2__60_carry__1_i_7__0_n_0;
  wire PSUM2__60_carry__1_i_7__1_n_0;
  wire PSUM2__60_carry__1_i_7__2_n_0;
  wire PSUM2__60_carry__1_i_7_n_0;
  wire PSUM2__60_carry__1_i_8__0_n_0;
  wire PSUM2__60_carry__1_i_8__1_n_0;
  wire PSUM2__60_carry__1_i_8__2_n_0;
  wire PSUM2__60_carry__1_i_8_n_0;
  wire PSUM2__60_carry__1_i_9__0_n_0;
  wire PSUM2__60_carry__1_i_9__1_n_0;
  wire PSUM2__60_carry__1_i_9__2_n_0;
  wire PSUM2__60_carry__1_i_9_n_0;
  wire PSUM2__60_carry__2_i_1__0_n_0;
  wire PSUM2__60_carry__2_i_1__1_n_0;
  wire PSUM2__60_carry__2_i_1__2_n_0;
  wire PSUM2__60_carry__2_i_1_n_0;
  wire PSUM2__60_carry_i_1__0_n_0;
  wire PSUM2__60_carry_i_1__1_n_0;
  wire PSUM2__60_carry_i_1__2_n_0;
  wire PSUM2__60_carry_i_1_n_0;
  wire PSUM2__60_carry_i_2__0_n_0;
  wire PSUM2__60_carry_i_2__1_n_0;
  wire PSUM2__60_carry_i_2__2_n_0;
  wire PSUM2__60_carry_i_2_n_0;
  wire PSUM2__60_carry_i_3__0_n_0;
  wire PSUM2__60_carry_i_3__1_n_0;
  wire PSUM2__60_carry_i_3__2_n_0;
  wire PSUM2__60_carry_i_3_n_0;
  wire PSUM2__60_carry_i_4__0_n_0;
  wire PSUM2__60_carry_i_4__1_n_0;
  wire PSUM2__60_carry_i_4__2_n_0;
  wire PSUM2__60_carry_i_4_n_0;
  wire PSUM2__60_carry_i_5__0_n_0;
  wire PSUM2__60_carry_i_5__1_n_0;
  wire PSUM2__60_carry_i_5__2_n_0;
  wire PSUM2__60_carry_i_5_n_0;
  wire PSUM3__0_carry__0_i_10__0_n_0;
  wire PSUM3__0_carry__0_i_10__1_n_0;
  wire PSUM3__0_carry__0_i_10__2_n_0;
  wire PSUM3__0_carry__0_i_10_n_0;
  wire PSUM3__0_carry__0_i_11__0_n_0;
  wire PSUM3__0_carry__0_i_11__1_n_0;
  wire PSUM3__0_carry__0_i_11__2_n_0;
  wire PSUM3__0_carry__0_i_11_n_0;
  wire PSUM3__0_carry__0_i_12__0_n_0;
  wire PSUM3__0_carry__0_i_12__1_n_0;
  wire PSUM3__0_carry__0_i_12__2_n_0;
  wire PSUM3__0_carry__0_i_12_n_0;
  wire PSUM3__0_carry__0_i_13_n_0;
  wire PSUM3__0_carry__0_i_1__0_n_0;
  wire PSUM3__0_carry__0_i_1__1_n_0;
  wire PSUM3__0_carry__0_i_1__2_n_0;
  wire PSUM3__0_carry__0_i_1_n_0;
  wire PSUM3__0_carry__0_i_2__0_n_0;
  wire PSUM3__0_carry__0_i_2__1_n_0;
  wire PSUM3__0_carry__0_i_2__2_n_0;
  wire PSUM3__0_carry__0_i_2_n_0;
  wire PSUM3__0_carry__0_i_3__0_n_0;
  wire PSUM3__0_carry__0_i_3__1_n_0;
  wire PSUM3__0_carry__0_i_3__2_n_0;
  wire PSUM3__0_carry__0_i_3_n_0;
  wire PSUM3__0_carry__0_i_4__0_n_0;
  wire PSUM3__0_carry__0_i_4__1_n_0;
  wire PSUM3__0_carry__0_i_4__2_n_0;
  wire PSUM3__0_carry__0_i_4_n_0;
  wire PSUM3__0_carry__0_i_5__0_n_0;
  wire PSUM3__0_carry__0_i_5__1_n_0;
  wire PSUM3__0_carry__0_i_5__2_n_0;
  wire PSUM3__0_carry__0_i_5_n_0;
  wire PSUM3__0_carry__0_i_6__0_n_0;
  wire PSUM3__0_carry__0_i_6__1_n_0;
  wire PSUM3__0_carry__0_i_6__2_n_0;
  wire PSUM3__0_carry__0_i_6_n_0;
  wire PSUM3__0_carry__0_i_7__0_n_0;
  wire PSUM3__0_carry__0_i_7__1_n_0;
  wire PSUM3__0_carry__0_i_7__2_n_0;
  wire PSUM3__0_carry__0_i_7_n_0;
  wire PSUM3__0_carry__0_i_8__0_n_0;
  wire PSUM3__0_carry__0_i_8__1_n_0;
  wire PSUM3__0_carry__0_i_8__2_n_0;
  wire PSUM3__0_carry__0_i_8_n_0;
  wire PSUM3__0_carry__0_i_9__0_n_0;
  wire PSUM3__0_carry__0_i_9__1_n_0;
  wire PSUM3__0_carry__0_i_9__2_n_0;
  wire PSUM3__0_carry__0_i_9_n_0;
  wire PSUM3__0_carry__1_i_1__0_n_0;
  wire PSUM3__0_carry__1_i_1__1_n_0;
  wire PSUM3__0_carry__1_i_1__2_n_0;
  wire PSUM3__0_carry__1_i_1_n_0;
  wire PSUM3__0_carry__1_i_2__0_n_0;
  wire PSUM3__0_carry__1_i_2__1_n_0;
  wire PSUM3__0_carry__1_i_2__2_n_0;
  wire PSUM3__0_carry__1_i_2_n_0;
  wire PSUM3__0_carry__1_i_3__0_n_0;
  wire PSUM3__0_carry__1_i_3__1_n_0;
  wire PSUM3__0_carry__1_i_3__2_n_0;
  wire PSUM3__0_carry__1_i_3_n_0;
  wire PSUM3__0_carry__1_i_4__0_n_0;
  wire PSUM3__0_carry__1_i_4__1_n_0;
  wire PSUM3__0_carry__1_i_4__2_n_0;
  wire PSUM3__0_carry__1_i_4_n_0;
  wire PSUM3__0_carry_i_1__0_n_0;
  wire PSUM3__0_carry_i_1__1_n_0;
  wire PSUM3__0_carry_i_1__2_n_0;
  wire PSUM3__0_carry_i_1_n_0;
  wire PSUM3__0_carry_i_2__0_n_0;
  wire PSUM3__0_carry_i_2__1_n_0;
  wire PSUM3__0_carry_i_2__2_n_0;
  wire PSUM3__0_carry_i_2_n_0;
  wire PSUM3__0_carry_i_3__0_n_0;
  wire PSUM3__0_carry_i_3__1_n_0;
  wire PSUM3__0_carry_i_3__2_n_0;
  wire PSUM3__0_carry_i_3_n_0;
  wire PSUM3__0_carry_i_4__0_n_0;
  wire PSUM3__0_carry_i_4__1_n_0;
  wire PSUM3__0_carry_i_4__2_n_0;
  wire PSUM3__0_carry_i_4_n_0;
  wire PSUM3__0_carry_i_5__0_n_0;
  wire PSUM3__0_carry_i_5__1_n_0;
  wire PSUM3__0_carry_i_5__2_n_0;
  wire PSUM3__0_carry_i_5_n_0;
  wire PSUM3__0_carry_i_6__0_n_0;
  wire PSUM3__0_carry_i_6__1_n_0;
  wire PSUM3__0_carry_i_6__2_n_0;
  wire PSUM3__0_carry_i_6_n_0;
  wire PSUM3__0_carry_i_7__0_n_0;
  wire PSUM3__0_carry_i_7__1_n_0;
  wire PSUM3__0_carry_i_7__2_n_0;
  wire PSUM3__0_carry_i_7_n_0;
  wire PSUM3__0_carry_i_8__0_n_0;
  wire PSUM3__0_carry_i_8__1_n_0;
  wire PSUM3__0_carry_i_8__2_n_0;
  wire PSUM3__0_carry_i_8_n_0;
  wire PSUM3__30_carry__0_i_10__0_n_0;
  wire PSUM3__30_carry__0_i_10__1_n_0;
  wire PSUM3__30_carry__0_i_10__2_n_0;
  wire PSUM3__30_carry__0_i_10_n_0;
  wire PSUM3__30_carry__0_i_11__0_n_0;
  wire PSUM3__30_carry__0_i_11__1_n_0;
  wire PSUM3__30_carry__0_i_11__2_n_0;
  wire PSUM3__30_carry__0_i_11_n_0;
  wire PSUM3__30_carry__0_i_12__0_n_0;
  wire PSUM3__30_carry__0_i_12__1_n_0;
  wire PSUM3__30_carry__0_i_12__2_n_0;
  wire PSUM3__30_carry__0_i_12_n_0;
  wire PSUM3__30_carry__0_i_1__0_n_0;
  wire PSUM3__30_carry__0_i_1__1_n_0;
  wire PSUM3__30_carry__0_i_1__2_n_0;
  wire PSUM3__30_carry__0_i_1_n_0;
  wire PSUM3__30_carry__0_i_2__0_n_0;
  wire PSUM3__30_carry__0_i_2__1_n_0;
  wire PSUM3__30_carry__0_i_2__2_n_0;
  wire PSUM3__30_carry__0_i_2_n_0;
  wire PSUM3__30_carry__0_i_3__0_n_0;
  wire PSUM3__30_carry__0_i_3__1_n_0;
  wire PSUM3__30_carry__0_i_3__2_n_0;
  wire PSUM3__30_carry__0_i_3_n_0;
  wire PSUM3__30_carry__0_i_4__0_n_0;
  wire PSUM3__30_carry__0_i_4__1_n_0;
  wire PSUM3__30_carry__0_i_4__2_n_0;
  wire PSUM3__30_carry__0_i_4_n_0;
  wire PSUM3__30_carry__0_i_5__0_n_0;
  wire PSUM3__30_carry__0_i_5__1_n_0;
  wire PSUM3__30_carry__0_i_5__2_n_0;
  wire PSUM3__30_carry__0_i_5_n_0;
  wire PSUM3__30_carry__0_i_6__0_n_0;
  wire PSUM3__30_carry__0_i_6__1_n_0;
  wire PSUM3__30_carry__0_i_6__2_n_0;
  wire PSUM3__30_carry__0_i_6_n_0;
  wire PSUM3__30_carry__0_i_7__0_n_0;
  wire PSUM3__30_carry__0_i_7__1_n_0;
  wire PSUM3__30_carry__0_i_7__2_n_0;
  wire PSUM3__30_carry__0_i_7_n_0;
  wire PSUM3__30_carry__0_i_8__0_n_0;
  wire PSUM3__30_carry__0_i_8__1_n_0;
  wire PSUM3__30_carry__0_i_8__2_n_0;
  wire PSUM3__30_carry__0_i_8_n_0;
  wire PSUM3__30_carry__0_i_9__0_n_0;
  wire PSUM3__30_carry__0_i_9__1_n_0;
  wire PSUM3__30_carry__0_i_9__2_n_0;
  wire PSUM3__30_carry__0_i_9_n_0;
  wire PSUM3__30_carry__1_i_1__0_n_0;
  wire PSUM3__30_carry__1_i_1__1_n_0;
  wire PSUM3__30_carry__1_i_1__2_n_0;
  wire PSUM3__30_carry__1_i_1_n_0;
  wire PSUM3__30_carry__1_i_2__0_n_0;
  wire PSUM3__30_carry__1_i_2__1_n_0;
  wire PSUM3__30_carry__1_i_2__2_n_0;
  wire PSUM3__30_carry__1_i_2_n_0;
  wire PSUM3__30_carry__1_i_3__0_n_0;
  wire PSUM3__30_carry__1_i_3__1_n_0;
  wire PSUM3__30_carry__1_i_3__2_n_0;
  wire PSUM3__30_carry__1_i_3_n_0;
  wire PSUM3__30_carry__1_i_4__0_n_0;
  wire PSUM3__30_carry__1_i_4__1_n_0;
  wire PSUM3__30_carry__1_i_4__2_n_0;
  wire PSUM3__30_carry__1_i_4_n_0;
  wire PSUM3__30_carry_i_1__0_n_0;
  wire PSUM3__30_carry_i_1__1_n_0;
  wire PSUM3__30_carry_i_1__2_n_0;
  wire PSUM3__30_carry_i_1_n_0;
  wire PSUM3__30_carry_i_2__0_n_0;
  wire PSUM3__30_carry_i_2__1_n_0;
  wire PSUM3__30_carry_i_2__2_n_0;
  wire PSUM3__30_carry_i_2_n_0;
  wire PSUM3__30_carry_i_3__0_n_0;
  wire PSUM3__30_carry_i_3__1_n_0;
  wire PSUM3__30_carry_i_3__2_n_0;
  wire PSUM3__30_carry_i_3_n_0;
  wire PSUM3__30_carry_i_4__0_n_0;
  wire PSUM3__30_carry_i_4__1_n_0;
  wire PSUM3__30_carry_i_4__2_n_0;
  wire PSUM3__30_carry_i_4_n_0;
  wire PSUM3__30_carry_i_5__0_n_0;
  wire PSUM3__30_carry_i_5__1_n_0;
  wire PSUM3__30_carry_i_5__2_n_0;
  wire PSUM3__30_carry_i_5_n_0;
  wire PSUM3__30_carry_i_6__0_n_0;
  wire PSUM3__30_carry_i_6__1_n_0;
  wire PSUM3__30_carry_i_6__2_n_0;
  wire PSUM3__30_carry_i_6_n_0;
  wire PSUM3__30_carry_i_7__0_n_0;
  wire PSUM3__30_carry_i_7__1_n_0;
  wire PSUM3__30_carry_i_7__2_n_0;
  wire PSUM3__30_carry_i_7_n_0;
  wire PSUM3__30_carry_i_8__0_n_0;
  wire PSUM3__30_carry_i_8__1_n_0;
  wire PSUM3__30_carry_i_8__2_n_0;
  wire PSUM3__30_carry_i_8_n_0;
  wire PSUM3__60_carry__0_i_10__0_n_0;
  wire PSUM3__60_carry__0_i_10__1_n_0;
  wire PSUM3__60_carry__0_i_10__2_n_0;
  wire PSUM3__60_carry__0_i_10_n_0;
  wire PSUM3__60_carry__0_i_11__0_n_0;
  wire PSUM3__60_carry__0_i_11__1_n_0;
  wire PSUM3__60_carry__0_i_11__2_n_0;
  wire PSUM3__60_carry__0_i_11_n_0;
  wire PSUM3__60_carry__0_i_12__0_n_0;
  wire PSUM3__60_carry__0_i_12__1_n_0;
  wire PSUM3__60_carry__0_i_12__2_n_0;
  wire PSUM3__60_carry__0_i_12_n_0;
  wire PSUM3__60_carry__0_i_13__0_n_0;
  wire PSUM3__60_carry__0_i_13__1_n_0;
  wire PSUM3__60_carry__0_i_13__2_n_0;
  wire PSUM3__60_carry__0_i_13_n_0;
  wire PSUM3__60_carry__0_i_14__0_n_0;
  wire PSUM3__60_carry__0_i_14__1_n_0;
  wire PSUM3__60_carry__0_i_14__2_n_0;
  wire PSUM3__60_carry__0_i_14_n_0;
  wire PSUM3__60_carry__0_i_15__0_n_0;
  wire PSUM3__60_carry__0_i_15__1_n_0;
  wire PSUM3__60_carry__0_i_15__2_n_0;
  wire PSUM3__60_carry__0_i_15_n_0;
  wire PSUM3__60_carry__0_i_1__0_n_0;
  wire PSUM3__60_carry__0_i_1__1_n_0;
  wire PSUM3__60_carry__0_i_1__2_n_0;
  wire PSUM3__60_carry__0_i_1_n_0;
  wire PSUM3__60_carry__0_i_2__0_n_0;
  wire PSUM3__60_carry__0_i_2__1_n_0;
  wire PSUM3__60_carry__0_i_2__2_n_0;
  wire PSUM3__60_carry__0_i_2_n_0;
  wire PSUM3__60_carry__0_i_3__0_n_0;
  wire PSUM3__60_carry__0_i_3__1_n_0;
  wire PSUM3__60_carry__0_i_3__2_n_0;
  wire PSUM3__60_carry__0_i_3_n_0;
  wire PSUM3__60_carry__0_i_4__0_n_0;
  wire PSUM3__60_carry__0_i_4__1_n_0;
  wire PSUM3__60_carry__0_i_4__2_n_0;
  wire PSUM3__60_carry__0_i_4_n_0;
  wire PSUM3__60_carry__0_i_5__0_n_0;
  wire PSUM3__60_carry__0_i_5__1_n_0;
  wire PSUM3__60_carry__0_i_5__2_n_0;
  wire PSUM3__60_carry__0_i_5_n_0;
  wire PSUM3__60_carry__0_i_6__0_n_0;
  wire PSUM3__60_carry__0_i_6__1_n_0;
  wire PSUM3__60_carry__0_i_6__2_n_0;
  wire PSUM3__60_carry__0_i_6_n_0;
  wire PSUM3__60_carry__0_i_7__0_n_0;
  wire PSUM3__60_carry__0_i_7__1_n_0;
  wire PSUM3__60_carry__0_i_7__2_n_0;
  wire PSUM3__60_carry__0_i_7_n_0;
  wire PSUM3__60_carry__0_i_8__0_n_0;
  wire PSUM3__60_carry__0_i_8__1_n_0;
  wire PSUM3__60_carry__0_i_8__2_n_0;
  wire PSUM3__60_carry__0_i_8_n_0;
  wire PSUM3__60_carry__0_i_9__0_n_0;
  wire PSUM3__60_carry__0_i_9__1_n_0;
  wire PSUM3__60_carry__0_i_9__2_n_0;
  wire PSUM3__60_carry__0_i_9_n_0;
  wire PSUM3__60_carry__1_i_10__0_n_0;
  wire PSUM3__60_carry__1_i_10__1_n_0;
  wire PSUM3__60_carry__1_i_10__2_n_0;
  wire PSUM3__60_carry__1_i_10_n_0;
  wire PSUM3__60_carry__1_i_11__0_n_0;
  wire PSUM3__60_carry__1_i_11__1_n_0;
  wire PSUM3__60_carry__1_i_11__2_n_0;
  wire PSUM3__60_carry__1_i_11_n_0;
  wire PSUM3__60_carry__1_i_12__0_n_0;
  wire PSUM3__60_carry__1_i_12__1_n_0;
  wire PSUM3__60_carry__1_i_12__2_n_0;
  wire PSUM3__60_carry__1_i_12_n_0;
  wire PSUM3__60_carry__1_i_13__0_n_0;
  wire PSUM3__60_carry__1_i_13__1_n_0;
  wire PSUM3__60_carry__1_i_13__2_n_0;
  wire PSUM3__60_carry__1_i_13_n_0;
  wire PSUM3__60_carry__1_i_14__0_n_0;
  wire PSUM3__60_carry__1_i_14__1_n_0;
  wire PSUM3__60_carry__1_i_14__2_n_0;
  wire PSUM3__60_carry__1_i_14_n_0;
  wire PSUM3__60_carry__1_i_15__0_n_0;
  wire PSUM3__60_carry__1_i_15__1_n_0;
  wire PSUM3__60_carry__1_i_15__2_n_0;
  wire PSUM3__60_carry__1_i_15_n_0;
  wire PSUM3__60_carry__1_i_1__0_n_0;
  wire PSUM3__60_carry__1_i_1__1_n_0;
  wire PSUM3__60_carry__1_i_1__2_n_0;
  wire PSUM3__60_carry__1_i_1_n_0;
  wire PSUM3__60_carry__1_i_2__0_n_0;
  wire PSUM3__60_carry__1_i_2__1_n_0;
  wire PSUM3__60_carry__1_i_2__2_n_0;
  wire PSUM3__60_carry__1_i_2_n_0;
  wire PSUM3__60_carry__1_i_3__0_n_0;
  wire PSUM3__60_carry__1_i_3__1_n_0;
  wire PSUM3__60_carry__1_i_3__2_n_0;
  wire PSUM3__60_carry__1_i_3_n_0;
  wire PSUM3__60_carry__1_i_4__0_n_0;
  wire PSUM3__60_carry__1_i_4__1_n_0;
  wire PSUM3__60_carry__1_i_4__2_n_0;
  wire PSUM3__60_carry__1_i_4_n_0;
  wire PSUM3__60_carry__1_i_5__0_n_0;
  wire PSUM3__60_carry__1_i_5__1_n_0;
  wire PSUM3__60_carry__1_i_5__2_n_0;
  wire PSUM3__60_carry__1_i_5_n_0;
  wire PSUM3__60_carry__1_i_6__0_n_0;
  wire PSUM3__60_carry__1_i_6__1_n_0;
  wire PSUM3__60_carry__1_i_6__2_n_0;
  wire PSUM3__60_carry__1_i_6_n_0;
  wire PSUM3__60_carry__1_i_7__0_n_0;
  wire PSUM3__60_carry__1_i_7__1_n_0;
  wire PSUM3__60_carry__1_i_7__2_n_0;
  wire PSUM3__60_carry__1_i_7_n_0;
  wire PSUM3__60_carry__1_i_8__0_n_0;
  wire PSUM3__60_carry__1_i_8__1_n_0;
  wire PSUM3__60_carry__1_i_8__2_n_0;
  wire PSUM3__60_carry__1_i_8_n_0;
  wire PSUM3__60_carry__1_i_9__0_n_0;
  wire PSUM3__60_carry__1_i_9__1_n_0;
  wire PSUM3__60_carry__1_i_9__2_n_0;
  wire PSUM3__60_carry__1_i_9_n_0;
  wire PSUM3__60_carry__2_i_1__0_n_0;
  wire PSUM3__60_carry__2_i_1__1_n_0;
  wire PSUM3__60_carry__2_i_1__2_n_0;
  wire PSUM3__60_carry__2_i_1_n_0;
  wire PSUM3__60_carry_i_1__0_n_0;
  wire PSUM3__60_carry_i_1__1_n_0;
  wire PSUM3__60_carry_i_1__2_n_0;
  wire PSUM3__60_carry_i_1_n_0;
  wire PSUM3__60_carry_i_2__0_n_0;
  wire PSUM3__60_carry_i_2__1_n_0;
  wire PSUM3__60_carry_i_2__2_n_0;
  wire PSUM3__60_carry_i_2_n_0;
  wire PSUM3__60_carry_i_3__0_n_0;
  wire PSUM3__60_carry_i_3__1_n_0;
  wire PSUM3__60_carry_i_3__2_n_0;
  wire PSUM3__60_carry_i_3_n_0;
  wire PSUM3__60_carry_i_4__0_n_0;
  wire PSUM3__60_carry_i_4__1_n_0;
  wire PSUM3__60_carry_i_4__2_n_0;
  wire PSUM3__60_carry_i_4_n_0;
  wire PSUM3__60_carry_i_5__0_n_0;
  wire PSUM3__60_carry_i_5__1_n_0;
  wire PSUM3__60_carry_i_5__2_n_0;
  wire PSUM3__60_carry_i_5_n_0;
  wire PSUM3_i_25_n_0;
  wire PSUM3_i_26_n_0;
  wire \Q[0]_i_1__4_n_0 ;
  wire \Q[0]_i_3_n_0 ;
  wire \Q[109]_i_2_n_0 ;
  wire \Q[109]_i_3_n_0 ;
  wire \Q[10]_i_2__0_n_0 ;
  wire \Q[10]_i_2__1_n_0 ;
  wire \Q[10]_i_2_n_0 ;
  wire \Q[10]_i_3__0_n_0 ;
  wire \Q[10]_i_3__1_n_0 ;
  wire \Q[10]_i_3_n_0 ;
  wire \Q[10]_i_4__0_n_0 ;
  wire \Q[10]_i_4_n_0 ;
  wire \Q[10]_i_5_n_0 ;
  wire \Q[10]_i_6_n_0 ;
  wire \Q[10]_i_7_n_0 ;
  wire \Q[112]_i_2_n_0 ;
  wire \Q[11]_i_10_n_0 ;
  wire \Q[11]_i_11_n_0 ;
  wire \Q[11]_i_16_n_0 ;
  wire \Q[11]_i_17_n_0 ;
  wire \Q[11]_i_2__0_n_0 ;
  wire \Q[11]_i_2__1_n_0 ;
  wire \Q[11]_i_2_n_0 ;
  wire \Q[11]_i_3__0_n_0 ;
  wire \Q[11]_i_3__1_n_0 ;
  wire \Q[11]_i_3_n_0 ;
  wire \Q[11]_i_4__0_n_0 ;
  wire \Q[11]_i_4__1_n_0 ;
  wire \Q[11]_i_4_n_0 ;
  wire \Q[11]_i_5__0_n_0 ;
  wire \Q[11]_i_5__1_n_0 ;
  wire \Q[11]_i_5_n_0 ;
  wire \Q[11]_i_6__0_n_0 ;
  wire \Q[11]_i_6_n_0 ;
  wire \Q[11]_i_7__0_n_0 ;
  wire \Q[11]_i_7_n_0 ;
  wire \Q[11]_i_9_n_0 ;
  wire \Q[123]_i_3_n_0 ;
  wire \Q[123]_i_5_n_0 ;
  wire \Q[123]_i_6_n_0 ;
  wire \Q[124]_i_3_n_0 ;
  wire \Q[125]_i_2_n_0 ;
  wire \Q[12]_i_10_n_0 ;
  wire \Q[12]_i_11__0_n_0 ;
  wire \Q[12]_i_11__1_n_0 ;
  wire \Q[12]_i_11_n_0 ;
  wire \Q[12]_i_12__0_n_0 ;
  wire \Q[12]_i_12__1_n_0 ;
  wire \Q[12]_i_12_n_0 ;
  wire \Q[12]_i_13__0_n_0 ;
  wire \Q[12]_i_13__1_n_0 ;
  wire \Q[12]_i_13_n_0 ;
  wire \Q[12]_i_14__0_n_0 ;
  wire \Q[12]_i_14_n_0 ;
  wire \Q[12]_i_15__0_n_0 ;
  wire \Q[12]_i_15_n_0 ;
  wire \Q[12]_i_16__0_n_0 ;
  wire \Q[12]_i_16_n_0 ;
  wire \Q[12]_i_17__0_n_0 ;
  wire \Q[12]_i_17_n_0 ;
  wire \Q[12]_i_18__0_n_0 ;
  wire \Q[12]_i_18_n_0 ;
  wire \Q[12]_i_19__0_n_0 ;
  wire \Q[12]_i_19_n_0 ;
  wire \Q[12]_i_20_n_0 ;
  wire \Q[12]_i_21_n_0 ;
  wire \Q[12]_i_22_n_0 ;
  wire \Q[12]_i_2__0_n_0 ;
  wire \Q[12]_i_2__1_n_0 ;
  wire \Q[12]_i_2_n_0 ;
  wire \Q[12]_i_3__0_n_0 ;
  wire \Q[12]_i_3__1_n_0 ;
  wire \Q[12]_i_3__2_n_0 ;
  wire \Q[12]_i_3__3_n_0 ;
  wire \Q[12]_i_4__0_n_0 ;
  wire \Q[12]_i_4__1_n_0 ;
  wire \Q[12]_i_4__2_n_0 ;
  wire \Q[12]_i_5__0_n_0 ;
  wire \Q[12]_i_5__1_n_0 ;
  wire \Q[12]_i_5__2_n_0 ;
  wire \Q[12]_i_6__0_n_0 ;
  wire \Q[12]_i_6__1_n_0 ;
  wire \Q[12]_i_7__0_n_0 ;
  wire \Q[12]_i_7_n_0 ;
  wire \Q[12]_i_8__0_n_0 ;
  wire \Q[12]_i_8_n_0 ;
  wire \Q[12]_i_9__0_n_0 ;
  wire \Q[12]_i_9_n_0 ;
  wire \Q[13]_i_10_n_0 ;
  wire \Q[13]_i_11_n_0 ;
  wire \Q[13]_i_12_n_0 ;
  wire \Q[13]_i_13_n_0 ;
  wire \Q[13]_i_14_n_0 ;
  wire \Q[13]_i_15_n_0 ;
  wire \Q[13]_i_16_n_0 ;
  wire \Q[13]_i_2__0_n_0 ;
  wire \Q[13]_i_2__1_n_0 ;
  wire \Q[13]_i_2_n_0 ;
  wire \Q[13]_i_3__0_n_0 ;
  wire \Q[13]_i_3_n_0 ;
  wire \Q[13]_i_4__0_n_0 ;
  wire \Q[13]_i_4_n_0 ;
  wire \Q[13]_i_5__0_n_0 ;
  wire \Q[13]_i_5_n_0 ;
  wire \Q[13]_i_6__0_n_0 ;
  wire \Q[13]_i_6_n_0 ;
  wire \Q[13]_i_7__0_n_0 ;
  wire \Q[13]_i_7_n_0 ;
  wire \Q[13]_i_8__0_n_0 ;
  wire \Q[13]_i_8_n_0 ;
  wire \Q[13]_i_9__0_n_0 ;
  wire \Q[13]_i_9_n_0 ;
  wire \Q[14]_i_2__0_n_0 ;
  wire \Q[14]_i_2__1_n_0 ;
  wire \Q[14]_i_2_n_0 ;
  wire \Q[14]_i_3__0_n_0 ;
  wire \Q[14]_i_3_n_0 ;
  wire \Q[14]_i_4__0_n_0 ;
  wire \Q[14]_i_4_n_0 ;
  wire \Q[14]_i_5_n_0 ;
  wire \Q[14]_i_6_n_0 ;
  wire \Q[14]_i_7_n_0 ;
  wire \Q[14]_i_8_n_0 ;
  wire \Q[14]_i_9_n_0 ;
  wire \Q[158]_rep__0_i_1_n_0 ;
  wire \Q[158]_rep__1_i_1_n_0 ;
  wire \Q[158]_rep__2_i_1_n_0 ;
  wire \Q[158]_rep__3_i_1_n_0 ;
  wire \Q[158]_rep__4_i_1_n_0 ;
  wire \Q[158]_rep_i_1_n_0 ;
  wire \Q[15]_i_10_n_0 ;
  wire \Q[15]_i_12_n_0 ;
  wire \Q[15]_i_13_n_0 ;
  wire \Q[15]_i_14_n_0 ;
  wire \Q[15]_i_15_n_0 ;
  wire \Q[15]_i_16_n_0 ;
  wire \Q[15]_i_17_n_0 ;
  wire \Q[15]_i_18_n_0 ;
  wire \Q[15]_i_19_n_0 ;
  wire \Q[15]_i_20_n_0 ;
  wire \Q[15]_i_21_n_0 ;
  wire \Q[15]_i_2__0_n_0 ;
  wire \Q[15]_i_2__1_n_0 ;
  wire \Q[15]_i_2__2_n_0 ;
  wire \Q[15]_i_2_n_0 ;
  wire \Q[15]_i_3__0_n_0 ;
  wire \Q[15]_i_3__1_n_0 ;
  wire \Q[15]_i_3_n_0 ;
  wire \Q[15]_i_4__0_n_0 ;
  wire \Q[15]_i_4_n_0 ;
  wire \Q[15]_i_5_n_0 ;
  wire \Q[15]_i_6__0_n_0 ;
  wire \Q[15]_i_6_n_0 ;
  wire \Q[15]_i_7__0_n_0 ;
  wire \Q[15]_i_7_n_0 ;
  wire \Q[15]_i_8_n_0 ;
  wire \Q[15]_i_9_n_0 ;
  wire \Q[160]_i_2_n_0 ;
  wire \Q[161]_i_2_n_0 ;
  wire \Q[161]_i_4_n_0 ;
  wire \Q[169]_i_2_n_0 ;
  wire \Q[16]_i_10__0_n_0 ;
  wire \Q[16]_i_10_n_0 ;
  wire \Q[16]_i_11__0_n_0 ;
  wire \Q[16]_i_11__1_n_0 ;
  wire \Q[16]_i_11_n_0 ;
  wire \Q[16]_i_12__0_n_0 ;
  wire \Q[16]_i_12__1_n_0 ;
  wire \Q[16]_i_12_n_0 ;
  wire \Q[16]_i_13__0_n_0 ;
  wire \Q[16]_i_13_n_0 ;
  wire \Q[16]_i_14__0_n_0 ;
  wire \Q[16]_i_14_n_0 ;
  wire \Q[16]_i_15__0_n_0 ;
  wire \Q[16]_i_15_n_0 ;
  wire \Q[16]_i_16__0_n_0 ;
  wire \Q[16]_i_16_n_0 ;
  wire \Q[16]_i_17_n_0 ;
  wire \Q[16]_i_18_n_0 ;
  wire \Q[16]_i_19_n_0 ;
  wire \Q[16]_i_20_n_0 ;
  wire \Q[16]_i_21_n_0 ;
  wire \Q[16]_i_22_n_0 ;
  wire \Q[16]_i_2__0_n_0 ;
  wire \Q[16]_i_2__1_n_0 ;
  wire \Q[16]_i_2__2_n_0 ;
  wire \Q[16]_i_2__3_n_0 ;
  wire \Q[16]_i_2_n_0 ;
  wire \Q[16]_i_3__0_n_0 ;
  wire \Q[16]_i_3__1_n_0 ;
  wire \Q[16]_i_3__2_n_0 ;
  wire \Q[16]_i_3__3_n_0 ;
  wire \Q[16]_i_4__0_n_0 ;
  wire \Q[16]_i_4__1_n_0 ;
  wire \Q[16]_i_4__2_n_0 ;
  wire \Q[16]_i_5__0_n_0 ;
  wire \Q[16]_i_5__1_n_0 ;
  wire \Q[16]_i_6__0_n_0 ;
  wire \Q[16]_i_7__0_n_0 ;
  wire \Q[16]_i_7_n_0 ;
  wire \Q[16]_i_8__0_n_0 ;
  wire \Q[16]_i_8_n_0 ;
  wire \Q[16]_i_9__0_n_0 ;
  wire \Q[16]_i_9_n_0 ;
  wire \Q[170]_rep__0_i_1_n_0 ;
  wire \Q[170]_rep__1_i_1_n_0 ;
  wire \Q[170]_rep__2_i_1_n_0 ;
  wire \Q[170]_rep__3_i_1_n_0 ;
  wire \Q[170]_rep_i_1_n_0 ;
  wire \Q[171]_i_100_n_0 ;
  wire \Q[171]_i_101_n_0 ;
  wire \Q[171]_i_102_n_0 ;
  wire \Q[171]_i_13_n_0 ;
  wire \Q[171]_i_14_n_0 ;
  wire \Q[171]_i_15_n_0 ;
  wire \Q[171]_i_17_n_0 ;
  wire \Q[171]_i_18_n_0 ;
  wire \Q[171]_i_19_n_0 ;
  wire \Q[171]_i_20_n_0 ;
  wire \Q[171]_i_21_n_0 ;
  wire \Q[171]_i_22_n_0 ;
  wire \Q[171]_i_23_n_0 ;
  wire \Q[171]_i_24_n_0 ;
  wire \Q[171]_i_26_n_0 ;
  wire \Q[171]_i_27_n_0 ;
  wire \Q[171]_i_28_n_0 ;
  wire \Q[171]_i_29_n_0 ;
  wire \Q[171]_i_2_n_0 ;
  wire \Q[171]_i_30_n_0 ;
  wire \Q[171]_i_31_n_0 ;
  wire \Q[171]_i_32_n_0 ;
  wire \Q[171]_i_33_n_0 ;
  wire \Q[171]_i_35_n_0 ;
  wire \Q[171]_i_36_n_0 ;
  wire \Q[171]_i_37_n_0 ;
  wire \Q[171]_i_38_n_0 ;
  wire \Q[171]_i_40_n_0 ;
  wire \Q[171]_i_41_n_0 ;
  wire \Q[171]_i_42_n_0 ;
  wire \Q[171]_i_43_n_0 ;
  wire \Q[171]_i_44_n_0 ;
  wire \Q[171]_i_45_n_0 ;
  wire \Q[171]_i_46_n_0 ;
  wire \Q[171]_i_47_n_0 ;
  wire \Q[171]_i_49_n_0 ;
  wire \Q[171]_i_4_n_0 ;
  wire \Q[171]_i_50_n_0 ;
  wire \Q[171]_i_51_n_0 ;
  wire \Q[171]_i_52_n_0 ;
  wire \Q[171]_i_53_n_0 ;
  wire \Q[171]_i_54_n_0 ;
  wire \Q[171]_i_55_n_0 ;
  wire \Q[171]_i_56_n_0 ;
  wire \Q[171]_i_57_n_0 ;
  wire \Q[171]_i_58_n_0 ;
  wire \Q[171]_i_59_n_0 ;
  wire \Q[171]_i_5_n_0 ;
  wire \Q[171]_i_60_n_0 ;
  wire \Q[171]_i_61_n_0 ;
  wire \Q[171]_i_62_n_0 ;
  wire \Q[171]_i_64_n_0 ;
  wire \Q[171]_i_65_n_0 ;
  wire \Q[171]_i_66_n_0 ;
  wire \Q[171]_i_67_n_0 ;
  wire \Q[171]_i_68_n_0 ;
  wire \Q[171]_i_69_n_0 ;
  wire \Q[171]_i_70_n_0 ;
  wire \Q[171]_i_71_n_0 ;
  wire \Q[171]_i_72_n_0 ;
  wire \Q[171]_i_74_n_0 ;
  wire \Q[171]_i_75_n_0 ;
  wire \Q[171]_i_76_n_0 ;
  wire \Q[171]_i_77_n_0 ;
  wire \Q[171]_i_78_n_0 ;
  wire \Q[171]_i_79_n_0 ;
  wire \Q[171]_i_7_n_0 ;
  wire \Q[171]_i_80_n_0 ;
  wire \Q[171]_i_81_n_0 ;
  wire \Q[171]_i_82_n_0 ;
  wire \Q[171]_i_83_n_0 ;
  wire \Q[171]_i_84_n_0 ;
  wire \Q[171]_i_85_n_0 ;
  wire \Q[171]_i_86_n_0 ;
  wire \Q[171]_i_87_n_0 ;
  wire \Q[171]_i_88_n_0 ;
  wire \Q[171]_i_89_n_0 ;
  wire \Q[171]_i_90_n_0 ;
  wire \Q[171]_i_91_n_0 ;
  wire \Q[171]_i_92_n_0 ;
  wire \Q[171]_i_93_n_0 ;
  wire \Q[171]_i_94_n_0 ;
  wire \Q[171]_i_95_n_0 ;
  wire \Q[171]_i_96_n_0 ;
  wire \Q[171]_i_97_n_0 ;
  wire \Q[171]_i_98_n_0 ;
  wire \Q[171]_i_99_n_0 ;
  wire \Q[171]_i_9_n_0 ;
  wire \Q[17]_i_10__0_n_0 ;
  wire \Q[17]_i_10_n_0 ;
  wire \Q[17]_i_11__0_n_0 ;
  wire \Q[17]_i_11_n_0 ;
  wire \Q[17]_i_12__0_n_0 ;
  wire \Q[17]_i_12_n_0 ;
  wire \Q[17]_i_13__0_n_0 ;
  wire \Q[17]_i_13_n_0 ;
  wire \Q[17]_i_14_n_0 ;
  wire \Q[17]_i_15_n_0 ;
  wire \Q[17]_i_16_n_0 ;
  wire \Q[17]_i_17_n_0 ;
  wire \Q[17]_i_18_n_0 ;
  wire \Q[17]_i_19_n_0 ;
  wire \Q[17]_i_20_n_0 ;
  wire \Q[17]_i_21_n_0 ;
  wire \Q[17]_i_2__0_n_0 ;
  wire \Q[17]_i_2__1_n_0 ;
  wire \Q[17]_i_2__2_n_0 ;
  wire \Q[17]_i_2_n_0 ;
  wire \Q[17]_i_3__0_n_0 ;
  wire \Q[17]_i_3__1_n_0 ;
  wire \Q[17]_i_3_n_0 ;
  wire \Q[17]_i_4__0_n_0 ;
  wire \Q[17]_i_4_n_0 ;
  wire \Q[17]_i_5__0_n_0 ;
  wire \Q[17]_i_5_n_0 ;
  wire \Q[17]_i_6__0_n_0 ;
  wire \Q[17]_i_6_n_0 ;
  wire \Q[17]_i_7__0_n_0 ;
  wire \Q[17]_i_7_n_0 ;
  wire \Q[17]_i_8__0_n_0 ;
  wire \Q[17]_i_8_n_0 ;
  wire \Q[17]_i_9__0_n_0 ;
  wire \Q[17]_i_9_n_0 ;
  wire \Q[18]_i_10__0_n_0 ;
  wire \Q[18]_i_10_n_0 ;
  wire \Q[18]_i_11__0_n_0 ;
  wire \Q[18]_i_11_n_0 ;
  wire \Q[18]_i_12__0_n_0 ;
  wire \Q[18]_i_12_n_0 ;
  wire \Q[18]_i_13_n_0 ;
  wire \Q[18]_i_14_n_0 ;
  wire \Q[18]_i_15_n_0 ;
  wire \Q[18]_i_16_n_0 ;
  wire \Q[18]_i_17_n_0 ;
  wire \Q[18]_i_2__0_n_0 ;
  wire \Q[18]_i_2__1_n_0 ;
  wire \Q[18]_i_2__2_n_0 ;
  wire \Q[18]_i_2_n_0 ;
  wire \Q[18]_i_3__0_n_0 ;
  wire \Q[18]_i_3_n_0 ;
  wire \Q[18]_i_4__0_n_0 ;
  wire \Q[18]_i_4_n_0 ;
  wire \Q[18]_i_5__0_n_0 ;
  wire \Q[18]_i_5_n_0 ;
  wire \Q[18]_i_6__0_n_0 ;
  wire \Q[18]_i_6_n_0 ;
  wire \Q[18]_i_7__0_n_0 ;
  wire \Q[18]_i_7_n_0 ;
  wire \Q[18]_i_8__0_n_0 ;
  wire \Q[18]_i_8_n_0 ;
  wire \Q[18]_i_9__0_n_0 ;
  wire \Q[18]_i_9_n_0 ;
  wire \Q[19]_i_10_n_0 ;
  wire \Q[19]_i_11_n_0 ;
  wire \Q[19]_i_12_n_0 ;
  wire \Q[19]_i_13_n_0 ;
  wire \Q[19]_i_2__0_n_0 ;
  wire \Q[19]_i_2__1_n_0 ;
  wire \Q[19]_i_2__2_n_0 ;
  wire \Q[19]_i_2_n_0 ;
  wire \Q[19]_i_3__0_n_0 ;
  wire \Q[19]_i_3__1_n_0 ;
  wire \Q[19]_i_3_n_0 ;
  wire \Q[19]_i_4__0_n_0 ;
  wire \Q[19]_i_4_n_0 ;
  wire \Q[19]_i_5__0_n_0 ;
  wire \Q[19]_i_5_n_0 ;
  wire \Q[19]_i_6_n_0 ;
  wire \Q[19]_i_7__0_n_0 ;
  wire \Q[19]_i_7_n_0 ;
  wire \Q[19]_i_8_n_0 ;
  wire \Q[19]_i_9_n_0 ;
  wire \Q[1]_i_2_n_0 ;
  wire \Q[20]_i_10__0_n_0 ;
  wire \Q[20]_i_10_n_0 ;
  wire \Q[20]_i_11__0_n_0 ;
  wire \Q[20]_i_11__1_n_0 ;
  wire \Q[20]_i_11_n_0 ;
  wire \Q[20]_i_12__0_n_0 ;
  wire \Q[20]_i_12__1_n_0 ;
  wire \Q[20]_i_12_n_0 ;
  wire \Q[20]_i_13__0_n_0 ;
  wire \Q[20]_i_13__1_n_0 ;
  wire \Q[20]_i_13_n_0 ;
  wire \Q[20]_i_14__0_n_0 ;
  wire \Q[20]_i_14__1_n_0 ;
  wire \Q[20]_i_14_n_0 ;
  wire \Q[20]_i_15_n_0 ;
  wire \Q[20]_i_16_n_0 ;
  wire \Q[20]_i_17_n_0 ;
  wire \Q[20]_i_18_n_0 ;
  wire \Q[20]_i_19_n_0 ;
  wire \Q[20]_i_20_n_0 ;
  wire \Q[20]_i_21_n_0 ;
  wire \Q[20]_i_22_n_0 ;
  wire \Q[20]_i_2__0_n_0 ;
  wire \Q[20]_i_2__1_n_0 ;
  wire \Q[20]_i_2__2_n_0 ;
  wire \Q[20]_i_2__3_n_0 ;
  wire \Q[20]_i_2_n_0 ;
  wire \Q[20]_i_3__0_n_0 ;
  wire \Q[20]_i_3__1_n_0 ;
  wire \Q[20]_i_3__2_n_0 ;
  wire \Q[20]_i_3__4_n_0 ;
  wire \Q[20]_i_4__0_n_0 ;
  wire \Q[20]_i_4__1_n_0 ;
  wire \Q[20]_i_4__2_n_0 ;
  wire \Q[20]_i_4__3_n_0 ;
  wire \Q[20]_i_5__0_n_0 ;
  wire \Q[20]_i_5__2_n_0 ;
  wire \Q[20]_i_6__0_n_0 ;
  wire \Q[20]_i_7__0_n_0 ;
  wire \Q[20]_i_7_n_0 ;
  wire \Q[20]_i_8__0_n_0 ;
  wire \Q[20]_i_8_n_0 ;
  wire \Q[20]_i_9__0_n_0 ;
  wire \Q[20]_i_9_n_0 ;
  wire \Q[21]_i_10__0_n_0 ;
  wire \Q[21]_i_10_n_0 ;
  wire \Q[21]_i_11__0_n_0 ;
  wire \Q[21]_i_11_n_0 ;
  wire \Q[21]_i_12__0_n_0 ;
  wire \Q[21]_i_12_n_0 ;
  wire \Q[21]_i_13_n_0 ;
  wire \Q[21]_i_2__0_n_0 ;
  wire \Q[21]_i_2__1_n_0 ;
  wire \Q[21]_i_2__2_n_0 ;
  wire \Q[21]_i_2_n_0 ;
  wire \Q[21]_i_3__0_n_0 ;
  wire \Q[21]_i_3__1_n_0 ;
  wire \Q[21]_i_3_n_0 ;
  wire \Q[21]_i_4__0_n_0 ;
  wire \Q[21]_i_4_n_0 ;
  wire \Q[21]_i_5_n_0 ;
  wire \Q[21]_i_6__0_n_0 ;
  wire \Q[21]_i_6_n_0 ;
  wire \Q[21]_i_7__0_n_0 ;
  wire \Q[21]_i_7_n_0 ;
  wire \Q[21]_i_8__0_n_0 ;
  wire \Q[21]_i_8_n_0 ;
  wire \Q[21]_i_9__0_n_0 ;
  wire \Q[21]_i_9_n_0 ;
  wire \Q[22]_i_10__0_n_0 ;
  wire \Q[22]_i_10_n_0 ;
  wire \Q[22]_i_11_n_0 ;
  wire \Q[22]_i_12__0_n_0 ;
  wire \Q[22]_i_12_n_0 ;
  wire \Q[22]_i_13__0_n_0 ;
  wire \Q[22]_i_13_n_0 ;
  wire \Q[22]_i_14__0_n_0 ;
  wire \Q[22]_i_14_n_0 ;
  wire \Q[22]_i_15__0_n_0 ;
  wire \Q[22]_i_15_n_0 ;
  wire \Q[22]_i_16__0_n_0 ;
  wire \Q[22]_i_16_n_0 ;
  wire \Q[22]_i_17__0_n_0 ;
  wire \Q[22]_i_17_n_0 ;
  wire \Q[22]_i_18__0_n_0 ;
  wire \Q[22]_i_18_n_0 ;
  wire \Q[22]_i_2__0_n_0 ;
  wire \Q[22]_i_2_n_0 ;
  wire \Q[22]_i_3__0_n_0 ;
  wire \Q[22]_i_3_n_0 ;
  wire \Q[22]_i_4_n_0 ;
  wire \Q[22]_i_5__0_n_0 ;
  wire \Q[22]_i_5_n_0 ;
  wire \Q[22]_i_6__0_n_0 ;
  wire \Q[22]_i_6_n_0 ;
  wire \Q[22]_i_7__0_n_0 ;
  wire \Q[22]_i_7_n_0 ;
  wire \Q[22]_i_8__0_n_0 ;
  wire \Q[22]_i_8_n_0 ;
  wire \Q[22]_i_9__0_n_0 ;
  wire \Q[22]_i_9_n_0 ;
  wire \Q[23]_i_11_n_0 ;
  wire \Q[23]_i_12_n_0 ;
  wire \Q[23]_i_13__0_n_0 ;
  wire \Q[23]_i_13_n_0 ;
  wire \Q[23]_i_14__0_n_0 ;
  wire \Q[23]_i_14_n_0 ;
  wire \Q[23]_i_15__0_n_0 ;
  wire \Q[23]_i_15_n_0 ;
  wire \Q[23]_i_16__0_n_0 ;
  wire \Q[23]_i_16_n_0 ;
  wire \Q[23]_i_17__0_n_0 ;
  wire \Q[23]_i_17_n_0 ;
  wire \Q[23]_i_18_n_0 ;
  wire \Q[23]_i_19_n_0 ;
  wire \Q[23]_i_20_n_0 ;
  wire \Q[23]_i_21_n_0 ;
  wire \Q[23]_i_22_n_0 ;
  wire \Q[23]_i_23_n_0 ;
  wire \Q[23]_i_2__0_n_0 ;
  wire \Q[23]_i_2_n_0 ;
  wire \Q[23]_i_3__0_n_0 ;
  wire \Q[23]_i_6__0_n_0 ;
  wire \Q[23]_i_7__0_n_0 ;
  wire \Q[23]_i_7_n_0 ;
  wire \Q[24]_i_10_n_0 ;
  wire \Q[24]_i_11_n_0 ;
  wire \Q[24]_i_12_n_0 ;
  wire \Q[24]_i_13_n_0 ;
  wire \Q[24]_i_14_n_0 ;
  wire \Q[24]_i_15_n_0 ;
  wire \Q[24]_i_16_n_0 ;
  wire \Q[24]_i_17_n_0 ;
  wire \Q[24]_i_18_n_0 ;
  wire \Q[24]_i_19_n_0 ;
  wire \Q[24]_i_2__0_n_0 ;
  wire \Q[24]_i_2__1_n_0 ;
  wire \Q[24]_i_2_n_0 ;
  wire \Q[24]_i_3__0_n_0 ;
  wire \Q[24]_i_3__1_n_0 ;
  wire \Q[24]_i_4__0_n_0 ;
  wire \Q[24]_i_4__1_n_0 ;
  wire \Q[24]_i_4_n_0 ;
  wire \Q[24]_i_5__0_n_0 ;
  wire \Q[24]_i_5__1_n_0 ;
  wire \Q[24]_i_5_n_0 ;
  wire \Q[24]_i_6__0_n_0 ;
  wire \Q[24]_i_7__0_n_0 ;
  wire \Q[24]_i_7_n_0 ;
  wire \Q[24]_i_8__0_n_0 ;
  wire \Q[24]_i_8_n_0 ;
  wire \Q[24]_i_9__0_n_0 ;
  wire \Q[24]_i_9_n_0 ;
  wire \Q[25]_i_2__0_n_0 ;
  wire \Q[25]_i_2_n_0 ;
  wire \Q[25]_i_3_n_0 ;
  wire \Q[25]_i_4_n_0 ;
  wire \Q[25]_i_5_n_0 ;
  wire \Q[25]_i_6_n_0 ;
  wire \Q[25]_i_8_n_0 ;
  wire \Q[26]_i_10__0_n_0 ;
  wire \Q[26]_i_10_n_0 ;
  wire \Q[26]_i_11__0_n_0 ;
  wire \Q[26]_i_11_n_0 ;
  wire \Q[26]_i_12__0_n_0 ;
  wire \Q[26]_i_12_n_0 ;
  wire \Q[26]_i_13__0_n_0 ;
  wire \Q[26]_i_13_n_0 ;
  wire \Q[26]_i_14__0_n_0 ;
  wire \Q[26]_i_14_n_0 ;
  wire \Q[26]_i_15__0_n_0 ;
  wire \Q[26]_i_15_n_0 ;
  wire \Q[26]_i_16__0_n_0 ;
  wire \Q[26]_i_16_n_0 ;
  wire \Q[26]_i_17__0_n_0 ;
  wire \Q[26]_i_17_n_0 ;
  wire \Q[26]_i_18__0_n_0 ;
  wire \Q[26]_i_18_n_0 ;
  wire \Q[26]_i_19_n_0 ;
  wire \Q[26]_i_20_n_0 ;
  wire \Q[26]_i_21_n_0 ;
  wire \Q[26]_i_22_n_0 ;
  wire \Q[26]_i_23_n_0 ;
  wire \Q[26]_i_2__0_n_0 ;
  wire \Q[26]_i_2_n_0 ;
  wire \Q[26]_i_3__0_n_0 ;
  wire \Q[26]_i_4__0_n_0 ;
  wire \Q[26]_i_4_n_0 ;
  wire \Q[26]_i_5__0_n_0 ;
  wire \Q[26]_i_5_n_0 ;
  wire \Q[26]_i_6__0_n_0 ;
  wire \Q[26]_i_6_n_0 ;
  wire \Q[26]_i_7__0_n_0 ;
  wire \Q[26]_i_7_n_0 ;
  wire \Q[26]_i_8__0_n_0 ;
  wire \Q[26]_i_9__0_n_0 ;
  wire \Q[26]_i_9_n_0 ;
  wire \Q[27]_i_13_n_0 ;
  wire \Q[27]_i_14_n_0 ;
  wire \Q[27]_i_15_n_0 ;
  wire \Q[27]_i_16_n_0 ;
  wire \Q[27]_i_17_n_0 ;
  wire \Q[27]_i_18_n_0 ;
  wire \Q[27]_i_2__0_n_0 ;
  wire \Q[27]_i_2__1_n_0 ;
  wire \Q[27]_i_2_n_0 ;
  wire \Q[27]_i_3__0_n_0 ;
  wire \Q[27]_i_3_n_0 ;
  wire \Q[27]_i_6_n_0 ;
  wire \Q[27]_i_7_n_0 ;
  wire \Q[28]_i_10_n_0 ;
  wire \Q[28]_i_11_n_0 ;
  wire \Q[28]_i_12_n_0 ;
  wire \Q[28]_i_13_n_0 ;
  wire \Q[28]_i_14_n_0 ;
  wire \Q[28]_i_15_n_0 ;
  wire \Q[28]_i_16_n_0 ;
  wire \Q[28]_i_17_n_0 ;
  wire \Q[28]_i_18_n_0 ;
  wire \Q[28]_i_19_n_0 ;
  wire \Q[28]_i_20_n_0 ;
  wire \Q[28]_i_21_n_0 ;
  wire \Q[28]_i_22_n_0 ;
  wire \Q[28]_i_23_n_0 ;
  wire \Q[28]_i_24_n_0 ;
  wire \Q[28]_i_2__0_n_0 ;
  wire \Q[28]_i_2__1_n_0 ;
  wire \Q[28]_i_2_n_0 ;
  wire \Q[28]_i_3__0_n_0 ;
  wire \Q[28]_i_3_n_0 ;
  wire \Q[28]_i_4__0_n_0 ;
  wire \Q[28]_i_4_n_0 ;
  wire \Q[28]_i_5__0_n_0 ;
  wire \Q[28]_i_5_n_0 ;
  wire \Q[28]_i_6_n_0 ;
  wire \Q[28]_i_7_n_0 ;
  wire \Q[28]_i_8_n_0 ;
  wire \Q[28]_i_9_n_0 ;
  wire \Q[29]_i_10__0_n_0 ;
  wire \Q[29]_i_10_n_0 ;
  wire \Q[29]_i_11__0_n_0 ;
  wire \Q[29]_i_11_n_0 ;
  wire \Q[29]_i_12__0_n_0 ;
  wire \Q[29]_i_12_n_0 ;
  wire \Q[29]_i_13__0_n_0 ;
  wire \Q[29]_i_13_n_0 ;
  wire \Q[29]_i_14_n_0 ;
  wire \Q[29]_i_15__0_n_0 ;
  wire \Q[29]_i_15_n_0 ;
  wire \Q[29]_i_16__0_n_0 ;
  wire \Q[29]_i_16_n_0 ;
  wire \Q[29]_i_17__0_n_0 ;
  wire \Q[29]_i_18__0_n_0 ;
  wire \Q[29]_i_19__0_n_0 ;
  wire \Q[29]_i_19_n_0 ;
  wire \Q[29]_i_20_n_0 ;
  wire \Q[29]_i_21_n_0 ;
  wire \Q[29]_i_22_n_0 ;
  wire \Q[29]_i_23_n_0 ;
  wire \Q[29]_i_24_n_0 ;
  wire \Q[29]_i_25_n_0 ;
  wire \Q[29]_i_26_n_0 ;
  wire \Q[29]_i_2__0_n_0 ;
  wire \Q[29]_i_2__1_n_0 ;
  wire \Q[29]_i_2__2_n_0 ;
  wire \Q[29]_i_3__1_n_0 ;
  wire \Q[29]_i_3_n_0 ;
  wire \Q[29]_i_4__0_n_0 ;
  wire \Q[29]_i_4__1_n_0 ;
  wire \Q[29]_i_4_n_0 ;
  wire \Q[29]_i_5__0_n_0 ;
  wire \Q[29]_i_5_n_0 ;
  wire \Q[29]_i_6__0_n_0 ;
  wire \Q[29]_i_6_n_0 ;
  wire \Q[29]_i_7__0_n_0 ;
  wire \Q[29]_i_7_n_0 ;
  wire \Q[29]_i_8__0_n_0 ;
  wire \Q[29]_i_8_n_0 ;
  wire \Q[29]_i_9_n_0 ;
  wire \Q[2]_i_2_n_0 ;
  wire \Q[30]_i_10__0_n_0 ;
  wire \Q[30]_i_10_n_0 ;
  wire \Q[30]_i_11__0_n_0 ;
  wire \Q[30]_i_11_n_0 ;
  wire \Q[30]_i_12__0_n_0 ;
  wire \Q[30]_i_12_n_0 ;
  wire \Q[30]_i_13__0_n_0 ;
  wire \Q[30]_i_13_n_0 ;
  wire \Q[30]_i_14__0_n_0 ;
  wire \Q[30]_i_14_n_0 ;
  wire \Q[30]_i_15_n_0 ;
  wire \Q[30]_i_16_n_0 ;
  wire \Q[30]_i_17_n_0 ;
  wire \Q[30]_i_22_n_0 ;
  wire \Q[30]_i_2__0_n_0 ;
  wire \Q[30]_i_2__1_n_0 ;
  wire \Q[30]_i_2__2_n_0 ;
  wire \Q[30]_i_2_n_0 ;
  wire \Q[30]_i_3__0_n_0 ;
  wire \Q[30]_i_4__0_n_0 ;
  wire \Q[30]_i_4__1_n_0 ;
  wire \Q[30]_i_4_n_0 ;
  wire \Q[30]_i_5__0_n_0 ;
  wire \Q[30]_i_5_n_0 ;
  wire \Q[30]_i_6__0_n_0 ;
  wire \Q[30]_i_6_n_0 ;
  wire \Q[30]_i_7_n_0 ;
  wire \Q[30]_i_8__0_n_0 ;
  wire \Q[30]_i_8_n_0 ;
  wire \Q[30]_i_9__0_n_0 ;
  wire \Q[30]_i_9_n_0 ;
  wire \Q[31]_i_10__0_n_0 ;
  wire \Q[31]_i_10_n_0 ;
  wire \Q[31]_i_11__0_n_0 ;
  wire \Q[31]_i_11_n_0 ;
  wire \Q[31]_i_12__0_n_0 ;
  wire \Q[31]_i_12_n_0 ;
  wire \Q[31]_i_13__0_n_0 ;
  wire \Q[31]_i_13_n_0 ;
  wire \Q[31]_i_14__0_n_0 ;
  wire \Q[31]_i_14_n_0 ;
  wire \Q[31]_i_15_n_0 ;
  wire \Q[31]_i_2__0_n_0 ;
  wire \Q[31]_i_2__1_n_0 ;
  wire \Q[31]_i_2__2_n_0 ;
  wire \Q[31]_i_2__3_n_0 ;
  wire \Q[31]_i_2__4_n_0 ;
  wire \Q[31]_i_2_n_0 ;
  wire \Q[31]_i_3__0_n_0 ;
  wire \Q[31]_i_3__2_n_0 ;
  wire \Q[31]_i_3__3_n_0 ;
  wire \Q[31]_i_3_n_0 ;
  wire \Q[31]_i_4__0_n_0 ;
  wire \Q[31]_i_4__1_n_0 ;
  wire \Q[31]_i_4__2_n_0 ;
  wire \Q[31]_i_4_n_0 ;
  wire \Q[31]_i_5__0_n_0 ;
  wire \Q[31]_i_5_n_0 ;
  wire \Q[31]_i_6__0_n_0 ;
  wire \Q[31]_i_6_n_0 ;
  wire \Q[31]_i_7__0_n_0 ;
  wire \Q[31]_i_7_n_0 ;
  wire \Q[31]_i_8_n_0 ;
  wire \Q[31]_i_9_n_0 ;
  wire \Q[32]_i_2__0_n_0 ;
  wire \Q[32]_i_2_n_0 ;
  wire \Q[32]_i_3_n_0 ;
  wire \Q[32]_i_4_n_0 ;
  wire \Q[33]_i_2__0_n_0 ;
  wire \Q[33]_i_2_n_0 ;
  wire \Q[33]_i_3__0_n_0 ;
  wire \Q[33]_i_3_n_0 ;
  wire \Q[34]_i_2__0_n_0 ;
  wire \Q[34]_i_2_n_0 ;
  wire \Q[34]_i_3__0_n_0 ;
  wire \Q[34]_i_3_n_0 ;
  wire \Q[34]_i_4_n_0 ;
  wire \Q[34]_i_5_n_0 ;
  wire \Q[34]_i_6_n_0 ;
  wire \Q[35]_i_10_n_0 ;
  wire \Q[35]_i_11_n_0 ;
  wire \Q[35]_i_16_n_0 ;
  wire \Q[35]_i_17_n_0 ;
  wire \Q[35]_i_18_n_0 ;
  wire \Q[35]_i_19_n_0 ;
  wire \Q[35]_i_20_n_0 ;
  wire \Q[35]_i_21_n_0 ;
  wire \Q[35]_i_22_n_0 ;
  wire \Q[35]_i_23_n_0 ;
  wire \Q[35]_i_24_n_0 ;
  wire \Q[35]_i_25_n_0 ;
  wire \Q[35]_i_26_n_0 ;
  wire \Q[35]_i_27_n_0 ;
  wire \Q[35]_i_28_n_0 ;
  wire \Q[35]_i_29_n_0 ;
  wire \Q[35]_i_2__0_n_0 ;
  wire \Q[35]_i_2_n_0 ;
  wire \Q[35]_i_32_n_0 ;
  wire \Q[35]_i_35_n_0 ;
  wire \Q[35]_i_36_n_0 ;
  wire \Q[35]_i_37_n_0 ;
  wire \Q[35]_i_38_n_0 ;
  wire \Q[35]_i_39_n_0 ;
  wire \Q[35]_i_3__0_n_0 ;
  wire \Q[35]_i_3_n_0 ;
  wire \Q[35]_i_40_n_0 ;
  wire \Q[35]_i_41_n_0 ;
  wire \Q[35]_i_42_n_0 ;
  wire \Q[35]_i_48_n_0 ;
  wire \Q[35]_i_4_n_0 ;
  wire \Q[35]_i_7_n_0 ;
  wire \Q[35]_i_8_n_0 ;
  wire \Q[35]_i_9_n_0 ;
  wire \Q[36]_i_2__0_n_0 ;
  wire \Q[36]_i_2__1_n_0 ;
  wire \Q[36]_i_3__0_n_0 ;
  wire \Q[36]_i_3_n_0 ;
  wire \Q[36]_i_4__0_n_0 ;
  wire \Q[36]_i_4_n_0 ;
  wire \Q[37]_i_2_n_0 ;
  wire \Q[37]_i_3_n_0 ;
  wire \Q[38]_i_2_n_0 ;
  wire \Q[39]_i_2_n_0 ;
  wire \Q[3]_i_2_n_0 ;
  wire \Q[3]_i_3_n_0 ;
  wire \Q[40]_i_2_n_0 ;
  wire \Q[41]_i_2_n_0 ;
  wire \Q[42]_i_2_n_0 ;
  wire \Q[43]_i_2_n_0 ;
  wire \Q[44]_i_2_n_0 ;
  wire \Q[45]_i_2_n_0 ;
  wire \Q[46]_i_10_n_0 ;
  wire \Q[46]_i_11_n_0 ;
  wire \Q[46]_i_12_n_0 ;
  wire \Q[46]_i_13_n_0 ;
  wire \Q[46]_i_14_n_0 ;
  wire \Q[46]_i_15_n_0 ;
  wire \Q[46]_i_16_n_0 ;
  wire \Q[46]_i_17_n_0 ;
  wire \Q[46]_i_2_n_0 ;
  wire \Q[46]_i_3_n_0 ;
  wire \Q[46]_i_4_n_0 ;
  wire \Q[46]_i_7_n_0 ;
  wire \Q[47]_i_1_n_0 ;
  wire \Q[47]_i_2_n_0 ;
  wire \Q[47]_i_4_n_0 ;
  wire \Q[47]_i_5_n_0 ;
  wire \Q[47]_i_6_n_0 ;
  wire \Q[47]_i_7_n_0 ;
  wire \Q[47]_i_8_n_0 ;
  wire \Q[47]_i_9_n_0 ;
  wire \Q[48]_i_10_n_0 ;
  wire \Q[48]_i_11_n_0 ;
  wire \Q[48]_i_12_n_0 ;
  wire \Q[48]_i_1_n_0 ;
  wire \Q[48]_i_2_n_0 ;
  wire \Q[48]_i_4_n_0 ;
  wire \Q[48]_i_5_n_0 ;
  wire \Q[48]_i_6_n_0 ;
  wire \Q[48]_i_7_n_0 ;
  wire \Q[48]_i_8_n_0 ;
  wire \Q[48]_i_9_n_0 ;
  wire \Q[49]_i_10_n_0 ;
  wire \Q[49]_i_11_n_0 ;
  wire \Q[49]_i_12_n_0 ;
  wire \Q[49]_i_13_n_0 ;
  wire \Q[49]_i_14_n_0 ;
  wire \Q[49]_i_15_n_0 ;
  wire \Q[49]_i_16_n_0 ;
  wire \Q[49]_i_19_n_0 ;
  wire \Q[49]_i_1_n_0 ;
  wire \Q[49]_i_20_n_0 ;
  wire \Q[49]_i_22_n_0 ;
  wire \Q[49]_i_23_n_0 ;
  wire \Q[49]_i_2_n_0 ;
  wire \Q[49]_i_33_n_0 ;
  wire \Q[49]_i_34_n_0 ;
  wire \Q[49]_i_36_n_0 ;
  wire \Q[49]_i_48_n_0 ;
  wire \Q[49]_i_4_n_0 ;
  wire \Q[49]_i_5_n_0 ;
  wire \Q[49]_i_7_n_0 ;
  wire \Q[49]_i_8_n_0 ;
  wire \Q[49]_i_9_n_0 ;
  wire \Q[4]_i_11_n_0 ;
  wire \Q[4]_i_12_n_0 ;
  wire \Q[4]_i_13_n_0 ;
  wire \Q[4]_i_14_n_0 ;
  wire \Q[4]_i_15_n_0 ;
  wire \Q[4]_i_16_n_0 ;
  wire \Q[4]_i_17_n_0 ;
  wire \Q[4]_i_18_n_0 ;
  wire \Q[4]_i_19_n_0 ;
  wire \Q[4]_i_20_n_0 ;
  wire \Q[4]_i_21_n_0 ;
  wire \Q[4]_i_22_n_0 ;
  wire \Q[4]_i_23_n_0 ;
  wire \Q[4]_i_24_n_0 ;
  wire \Q[4]_i_25_n_0 ;
  wire \Q[4]_i_26_n_0 ;
  wire \Q[4]_i_27_n_0 ;
  wire \Q[4]_i_2_n_0 ;
  wire \Q[4]_i_3__0_n_0 ;
  wire \Q[4]_i_3__1_n_0 ;
  wire \Q[4]_i_4__0_n_0 ;
  wire \Q[4]_i_4__1_n_0 ;
  wire \Q[4]_i_5__0_n_0 ;
  wire \Q[4]_i_5__1_n_0 ;
  wire \Q[4]_i_6__0_n_0 ;
  wire \Q[4]_i_7_n_0 ;
  wire \Q[4]_i_8_n_0 ;
  wire \Q[4]_i_9_n_0 ;
  wire \Q[50]_i_1_n_0 ;
  wire \Q[50]_i_2_n_0 ;
  wire \Q[51]_i_1_n_0 ;
  wire \Q[51]_i_2_n_0 ;
  wire \Q[52]_i_10_n_0 ;
  wire \Q[52]_i_11_n_0 ;
  wire \Q[52]_i_12_n_0 ;
  wire \Q[52]_i_13_n_0 ;
  wire \Q[52]_i_1_n_0 ;
  wire \Q[52]_i_2_n_0 ;
  wire \Q[52]_i_4_n_0 ;
  wire \Q[52]_i_5_n_0 ;
  wire \Q[52]_i_6_n_0 ;
  wire \Q[52]_i_7_n_0 ;
  wire \Q[52]_i_8_n_0 ;
  wire \Q[52]_i_9_n_0 ;
  wire \Q[53]_i_1_n_0 ;
  wire \Q[53]_i_2_n_0 ;
  wire \Q[54]_i_1_n_0 ;
  wire \Q[54]_i_2_n_0 ;
  wire \Q[55]_i_1__0_n_0 ;
  wire \Q[55]_i_2_n_0 ;
  wire \Q[56]_i_1__0_n_0 ;
  wire \Q[56]_i_2_n_0 ;
  wire \Q[57]_i_1__0_n_0 ;
  wire \Q[57]_i_2_n_0 ;
  wire \Q[58]_i_1__0_n_0 ;
  wire \Q[58]_i_2_n_0 ;
  wire \Q[59]_i_1__0_n_0 ;
  wire \Q[59]_i_2_n_0 ;
  wire \Q[5]_i_10_n_0 ;
  wire \Q[5]_i_2__0_n_0 ;
  wire \Q[5]_i_2__1_n_0 ;
  wire \Q[5]_i_2__2_n_0 ;
  wire \Q[5]_i_2_n_0 ;
  wire \Q[5]_i_3__0_n_0 ;
  wire \Q[5]_i_3__1_n_0 ;
  wire \Q[5]_i_3_n_0 ;
  wire \Q[5]_i_4_n_0 ;
  wire \Q[5]_i_5_n_0 ;
  wire \Q[60]_i_1__0_n_0 ;
  wire \Q[60]_i_2_n_0 ;
  wire \Q[61]_i_1__0_n_0 ;
  wire \Q[61]_i_2_n_0 ;
  wire \Q[62]_i_1__0_n_0 ;
  wire \Q[62]_i_2_n_0 ;
  wire \Q[63]_i_1__1_n_0 ;
  wire \Q[63]_i_1_n_0 ;
  wire \Q[63]_i_2_n_0 ;
  wire \Q[64]_i_1__0_n_0 ;
  wire \Q[64]_i_2_n_0 ;
  wire \Q[65]_i_10_n_0 ;
  wire \Q[65]_i_11_n_0 ;
  wire \Q[65]_i_12_n_0 ;
  wire \Q[65]_i_13_n_0 ;
  wire \Q[65]_i_14_n_0 ;
  wire \Q[65]_i_15_n_0 ;
  wire \Q[65]_i_17_n_0 ;
  wire \Q[65]_i_18_n_0 ;
  wire \Q[65]_i_19_n_0 ;
  wire \Q[65]_i_1__0_n_0 ;
  wire \Q[65]_i_20_n_0 ;
  wire \Q[65]_i_21_n_0 ;
  wire \Q[65]_i_22_n_0 ;
  wire \Q[65]_i_23_n_0 ;
  wire \Q[65]_i_2_n_0 ;
  wire \Q[65]_i_4_n_0 ;
  wire \Q[65]_i_5_n_0 ;
  wire \Q[65]_i_7_n_0 ;
  wire \Q[65]_i_8_n_0 ;
  wire \Q[65]_i_9_n_0 ;
  wire \Q[66]_i_10_n_0 ;
  wire \Q[66]_i_11_n_0 ;
  wire \Q[66]_i_12_n_0 ;
  wire \Q[66]_i_13_n_0 ;
  wire \Q[66]_i_14_n_0 ;
  wire \Q[66]_i_15_n_0 ;
  wire \Q[66]_i_16_n_0 ;
  wire \Q[66]_i_17_n_0 ;
  wire \Q[66]_i_18_n_0 ;
  wire \Q[66]_i_19_n_0 ;
  wire \Q[66]_i_1__0_n_0 ;
  wire \Q[66]_i_20_n_0 ;
  wire \Q[66]_i_2_n_0 ;
  wire \Q[66]_i_4_n_0 ;
  wire \Q[66]_i_5_n_0 ;
  wire \Q[66]_i_6_n_0 ;
  wire \Q[66]_i_7_n_0 ;
  wire \Q[66]_i_8_n_0 ;
  wire \Q[66]_i_9_n_0 ;
  wire \Q[67]_i_10__0_n_0 ;
  wire \Q[67]_i_10_n_0 ;
  wire \Q[67]_i_11__0_n_0 ;
  wire \Q[67]_i_11_n_0 ;
  wire \Q[67]_i_12__0_n_0 ;
  wire \Q[67]_i_12_n_0 ;
  wire \Q[67]_i_13__0_n_0 ;
  wire \Q[67]_i_13_n_0 ;
  wire \Q[67]_i_14__0_n_0 ;
  wire \Q[67]_i_14_n_0 ;
  wire \Q[67]_i_15_n_0 ;
  wire \Q[67]_i_16_n_0 ;
  wire \Q[67]_i_17_n_0 ;
  wire \Q[67]_i_18_n_0 ;
  wire \Q[67]_i_19_n_0 ;
  wire \Q[67]_i_1__0_n_0 ;
  wire \Q[67]_i_20_n_0 ;
  wire \Q[67]_i_21_n_0 ;
  wire \Q[67]_i_2_n_0 ;
  wire \Q[67]_i_4_n_0 ;
  wire \Q[67]_i_5_n_0 ;
  wire \Q[67]_i_6_n_0 ;
  wire \Q[67]_i_7_n_0 ;
  wire \Q[67]_i_8_n_0 ;
  wire \Q[67]_i_9__0_n_0 ;
  wire \Q[67]_i_9_n_0 ;
  wire \Q[68]_i_1__0_n_0 ;
  wire \Q[68]_i_2_n_0 ;
  wire \Q[69]_i_10_n_0 ;
  wire \Q[69]_i_11_n_0 ;
  wire \Q[69]_i_12_n_0 ;
  wire \Q[69]_i_13_n_0 ;
  wire \Q[69]_i_14_n_0 ;
  wire \Q[69]_i_15_n_0 ;
  wire \Q[69]_i_16_n_0 ;
  wire \Q[69]_i_17_n_0 ;
  wire \Q[69]_i_18_n_0 ;
  wire \Q[69]_i_19_n_0 ;
  wire \Q[69]_i_1__0_n_0 ;
  wire \Q[69]_i_20_n_0 ;
  wire \Q[69]_i_21_n_0 ;
  wire \Q[69]_i_22_n_0 ;
  wire \Q[69]_i_23_n_0 ;
  wire \Q[69]_i_24_n_0 ;
  wire \Q[69]_i_25_n_0 ;
  wire \Q[69]_i_26_n_0 ;
  wire \Q[69]_i_27_n_0 ;
  wire \Q[69]_i_28_n_0 ;
  wire \Q[69]_i_29_n_0 ;
  wire \Q[69]_i_2_n_0 ;
  wire \Q[69]_i_30_n_0 ;
  wire \Q[69]_i_31_n_0 ;
  wire \Q[69]_i_32_n_0 ;
  wire \Q[69]_i_33_n_0 ;
  wire \Q[69]_i_34_n_0 ;
  wire \Q[69]_i_35_n_0 ;
  wire \Q[69]_i_4_n_0 ;
  wire \Q[69]_i_5_n_0 ;
  wire \Q[69]_i_6_n_0 ;
  wire \Q[69]_i_7_n_0 ;
  wire \Q[69]_i_9_n_0 ;
  wire \Q[6]_i_2__0_n_0 ;
  wire \Q[6]_i_2_n_0 ;
  wire \Q[6]_i_3__0_n_0 ;
  wire \Q[6]_i_3_n_0 ;
  wire \Q[6]_i_4_n_0 ;
  wire \Q[70]_i_1__0_n_0 ;
  wire \Q[70]_i_2_n_0 ;
  wire \Q[71]_i_10_n_0 ;
  wire \Q[71]_i_11_n_0 ;
  wire \Q[71]_i_1__0_n_0 ;
  wire \Q[71]_i_2_n_0 ;
  wire \Q[71]_i_8_n_0 ;
  wire \Q[71]_i_9_n_0 ;
  wire \Q[72]_i_1__0_n_0 ;
  wire \Q[72]_i_2_n_0 ;
  wire \Q[73]_i_1__0_n_0 ;
  wire \Q[73]_i_2_n_0 ;
  wire \Q[74]_i_1__0_n_0 ;
  wire \Q[74]_i_2_n_0 ;
  wire \Q[75]_i_10_n_0 ;
  wire \Q[75]_i_11_n_0 ;
  wire \Q[75]_i_1__0_n_0 ;
  wire \Q[75]_i_2_n_0 ;
  wire \Q[75]_i_8_n_0 ;
  wire \Q[75]_i_9_n_0 ;
  wire \Q[76]_i_1__0_n_0 ;
  wire \Q[76]_i_2_n_0 ;
  wire \Q[77]_i_1__0_n_0 ;
  wire \Q[77]_i_2_n_0 ;
  wire \Q[77]_i_3_n_0 ;
  wire \Q[77]_i_4_n_0 ;
  wire \Q[77]_i_5_n_0 ;
  wire \Q[77]_i_6_n_0 ;
  wire \Q[78]_i_10_n_0 ;
  wire \Q[78]_i_11_n_0 ;
  wire \Q[78]_i_12_n_0 ;
  wire \Q[78]_i_13_n_0 ;
  wire \Q[78]_i_14_n_0 ;
  wire \Q[78]_i_15_n_0 ;
  wire \Q[78]_i_16_n_0 ;
  wire \Q[78]_i_17_n_0 ;
  wire \Q[78]_i_1__0_n_0 ;
  wire \Q[78]_i_2_n_0 ;
  wire \Q[78]_i_3_n_0 ;
  wire \Q[78]_i_4_n_0 ;
  wire \Q[78]_i_9_n_0 ;
  wire \Q[79]_i_10_n_0 ;
  wire \Q[79]_i_11_n_0 ;
  wire \Q[79]_i_2_n_0 ;
  wire \Q[79]_i_3_n_0 ;
  wire \Q[79]_i_4_n_0 ;
  wire \Q[79]_i_8_n_0 ;
  wire \Q[79]_i_9_n_0 ;
  wire \Q[7]_i_2__0_n_0 ;
  wire \Q[7]_i_2_n_0 ;
  wire \Q[7]_i_3__0_n_0 ;
  wire \Q[7]_i_3_n_0 ;
  wire \Q[7]_i_4_n_0 ;
  wire \Q[7]_i_5_n_0 ;
  wire \Q[83]_i_10_n_0 ;
  wire \Q[83]_i_11_n_0 ;
  wire \Q[83]_i_2_n_0 ;
  wire \Q[83]_i_3_n_0 ;
  wire \Q[83]_i_8_n_0 ;
  wire \Q[83]_i_9_n_0 ;
  wire \Q[87]_i_10_n_0 ;
  wire \Q[87]_i_11_n_0 ;
  wire \Q[87]_i_12_n_0 ;
  wire \Q[87]_i_4_n_0 ;
  wire \Q[87]_i_8_n_0 ;
  wire \Q[87]_i_9_n_0 ;
  wire \Q[88]_i_3_n_0 ;
  wire \Q[88]_i_4_n_0 ;
  wire \Q[88]_i_5_n_0 ;
  wire \Q[8]_i_10__0_n_0 ;
  wire \Q[8]_i_10_n_0 ;
  wire \Q[8]_i_11_n_0 ;
  wire \Q[8]_i_12_n_0 ;
  wire \Q[8]_i_13_n_0 ;
  wire \Q[8]_i_14_n_0 ;
  wire \Q[8]_i_15_n_0 ;
  wire \Q[8]_i_16_n_0 ;
  wire \Q[8]_i_17_n_0 ;
  wire \Q[8]_i_18_n_0 ;
  wire \Q[8]_i_19_n_0 ;
  wire \Q[8]_i_20_n_0 ;
  wire \Q[8]_i_21_n_0 ;
  wire \Q[8]_i_22_n_0 ;
  wire \Q[8]_i_2__0_n_0 ;
  wire \Q[8]_i_2__1_n_0 ;
  wire \Q[8]_i_2_n_0 ;
  wire \Q[8]_i_3__0_n_0 ;
  wire \Q[8]_i_3__1_n_0 ;
  wire \Q[8]_i_3__2_n_0 ;
  wire \Q[8]_i_3__3_n_0 ;
  wire \Q[8]_i_4__1_n_0 ;
  wire \Q[8]_i_4__2_n_0 ;
  wire \Q[8]_i_4_n_0 ;
  wire \Q[8]_i_5__0_n_0 ;
  wire \Q[8]_i_5__1_n_0 ;
  wire \Q[8]_i_5__2_n_0 ;
  wire \Q[8]_i_6__0_n_0 ;
  wire \Q[8]_i_6__1_n_0 ;
  wire \Q[8]_i_7__0_n_0 ;
  wire \Q[8]_i_7_n_0 ;
  wire \Q[8]_i_8__0_n_0 ;
  wire \Q[8]_i_8_n_0 ;
  wire \Q[8]_i_9__0_n_0 ;
  wire \Q[8]_i_9_n_0 ;
  wire \Q[90]_i_2_n_0 ;
  wire \Q[90]_i_3_n_0 ;
  wire \Q[90]_i_4_n_0 ;
  wire \Q[90]_i_5_n_0 ;
  wire \Q[90]_i_6_n_0 ;
  wire \Q[92]_i_2_n_0 ;
  wire \Q[92]_i_3_n_0 ;
  wire \Q[98]_i_2_n_0 ;
  wire \Q[98]_i_3_n_0 ;
  wire \Q[98]_i_4_n_0 ;
  wire \Q[9]_i_10__0_n_0 ;
  wire \Q[9]_i_10_n_0 ;
  wire \Q[9]_i_11__0_n_0 ;
  wire \Q[9]_i_11_n_0 ;
  wire \Q[9]_i_12__0_n_0 ;
  wire \Q[9]_i_12_n_0 ;
  wire \Q[9]_i_13__0_n_0 ;
  wire \Q[9]_i_13_n_0 ;
  wire \Q[9]_i_14_n_0 ;
  wire \Q[9]_i_15_n_0 ;
  wire \Q[9]_i_16_n_0 ;
  wire \Q[9]_i_2__0_n_0 ;
  wire \Q[9]_i_2__1_n_0 ;
  wire \Q[9]_i_2_n_0 ;
  wire \Q[9]_i_3__0_n_0 ;
  wire \Q[9]_i_3__1_n_0 ;
  wire \Q[9]_i_3__2_n_0 ;
  wire \Q[9]_i_4__0_n_0 ;
  wire \Q[9]_i_4__1_n_0 ;
  wire \Q[9]_i_4_n_0 ;
  wire \Q[9]_i_5__0_n_0 ;
  wire \Q[9]_i_5_n_0 ;
  wire \Q[9]_i_6__0_n_0 ;
  wire \Q[9]_i_6__1_n_0 ;
  wire \Q[9]_i_7__0_n_0 ;
  wire \Q[9]_i_8__0_n_0 ;
  wire \Q[9]_i_8_n_0 ;
  wire \Q[9]_i_9__0_n_0 ;
  wire \Q[9]_i_9_n_0 ;
  wire \Q_reg[12]_i_10_n_0 ;
  wire \Q_reg[12]_i_10_n_1 ;
  wire \Q_reg[12]_i_10_n_2 ;
  wire \Q_reg[12]_i_10_n_3 ;
  wire \Q_reg[12]_i_1_n_0 ;
  wire \Q_reg[12]_i_1_n_1 ;
  wire \Q_reg[12]_i_1_n_2 ;
  wire \Q_reg[12]_i_1_n_3 ;
  wire \Q_reg[12]_i_2__0_n_0 ;
  wire \Q_reg[12]_i_2__0_n_1 ;
  wire \Q_reg[12]_i_2__0_n_2 ;
  wire \Q_reg[12]_i_2__0_n_3 ;
  wire \Q_reg[12]_i_2_n_0 ;
  wire \Q_reg[12]_i_2_n_1 ;
  wire \Q_reg[12]_i_2_n_2 ;
  wire \Q_reg[12]_i_2_n_3 ;
  wire \Q_reg[16]_i_13_n_0 ;
  wire \Q_reg[16]_i_13_n_1 ;
  wire \Q_reg[16]_i_13_n_2 ;
  wire \Q_reg[16]_i_13_n_3 ;
  wire \Q_reg[16]_i_13_n_4 ;
  wire \Q_reg[16]_i_13_n_5 ;
  wire \Q_reg[16]_i_13_n_6 ;
  wire \Q_reg[16]_i_13_n_7 ;
  wire \Q_reg[16]_i_1_n_0 ;
  wire \Q_reg[16]_i_1_n_1 ;
  wire \Q_reg[16]_i_1_n_2 ;
  wire \Q_reg[16]_i_1_n_3 ;
  wire \Q_reg[16]_i_2_n_0 ;
  wire \Q_reg[16]_i_2_n_1 ;
  wire \Q_reg[16]_i_2_n_2 ;
  wire \Q_reg[16]_i_2_n_3 ;
  wire \Q_reg[16]_i_5_n_0 ;
  wire \Q_reg[16]_i_5_n_1 ;
  wire \Q_reg[16]_i_5_n_2 ;
  wire \Q_reg[16]_i_5_n_3 ;
  wire \Q_reg[16]_i_6_n_0 ;
  wire \Q_reg[16]_i_6_n_1 ;
  wire \Q_reg[16]_i_6_n_2 ;
  wire \Q_reg[16]_i_6_n_3 ;
  wire \Q_reg[171]_i_10_n_1 ;
  wire \Q_reg[171]_i_10_n_2 ;
  wire \Q_reg[171]_i_10_n_3 ;
  wire \Q_reg[171]_i_11_n_0 ;
  wire \Q_reg[171]_i_11_n_1 ;
  wire \Q_reg[171]_i_11_n_2 ;
  wire \Q_reg[171]_i_11_n_3 ;
  wire \Q_reg[171]_i_12_n_0 ;
  wire \Q_reg[171]_i_12_n_1 ;
  wire \Q_reg[171]_i_12_n_2 ;
  wire \Q_reg[171]_i_12_n_3 ;
  wire \Q_reg[171]_i_16_n_0 ;
  wire \Q_reg[171]_i_16_n_1 ;
  wire \Q_reg[171]_i_16_n_2 ;
  wire \Q_reg[171]_i_16_n_3 ;
  wire \Q_reg[171]_i_25_n_0 ;
  wire \Q_reg[171]_i_25_n_1 ;
  wire \Q_reg[171]_i_25_n_2 ;
  wire \Q_reg[171]_i_25_n_3 ;
  wire \Q_reg[171]_i_34_n_0 ;
  wire \Q_reg[171]_i_34_n_1 ;
  wire \Q_reg[171]_i_34_n_2 ;
  wire \Q_reg[171]_i_34_n_3 ;
  wire \Q_reg[171]_i_39_n_0 ;
  wire \Q_reg[171]_i_39_n_1 ;
  wire \Q_reg[171]_i_39_n_2 ;
  wire \Q_reg[171]_i_39_n_3 ;
  wire \Q_reg[171]_i_48_n_0 ;
  wire \Q_reg[171]_i_48_n_1 ;
  wire \Q_reg[171]_i_48_n_2 ;
  wire \Q_reg[171]_i_48_n_3 ;
  wire \Q_reg[171]_i_63_n_0 ;
  wire \Q_reg[171]_i_63_n_1 ;
  wire \Q_reg[171]_i_63_n_2 ;
  wire \Q_reg[171]_i_63_n_3 ;
  wire \Q_reg[171]_i_73_n_0 ;
  wire \Q_reg[171]_i_73_n_1 ;
  wire \Q_reg[171]_i_73_n_2 ;
  wire \Q_reg[171]_i_73_n_3 ;
  wire \Q_reg[171]_i_8_n_2 ;
  wire \Q_reg[171]_i_8_n_3 ;
  wire \Q_reg[20]_i_1_n_0 ;
  wire \Q_reg[20]_i_1_n_1 ;
  wire \Q_reg[20]_i_1_n_2 ;
  wire \Q_reg[20]_i_1_n_3 ;
  wire \Q_reg[20]_i_2_n_0 ;
  wire \Q_reg[20]_i_2_n_1 ;
  wire \Q_reg[20]_i_2_n_2 ;
  wire \Q_reg[20]_i_2_n_3 ;
  wire \Q_reg[20]_i_6_n_0 ;
  wire \Q_reg[20]_i_6_n_1 ;
  wire \Q_reg[20]_i_6_n_2 ;
  wire \Q_reg[20]_i_6_n_3 ;
  wire \Q_reg[22]_i_2_n_3 ;
  wire \Q_reg[22]_i_4_n_0 ;
  wire \Q_reg[22]_i_4_n_1 ;
  wire \Q_reg[22]_i_4_n_2 ;
  wire \Q_reg[22]_i_4_n_3 ;
  wire \Q_reg[23]_i_2_n_0 ;
  wire \Q_reg[23]_i_2_n_1 ;
  wire \Q_reg[23]_i_2_n_2 ;
  wire \Q_reg[23]_i_2_n_3 ;
  wire \Q_reg[24]_i_1_n_0 ;
  wire \Q_reg[24]_i_1_n_1 ;
  wire \Q_reg[24]_i_1_n_2 ;
  wire \Q_reg[24]_i_1_n_3 ;
  wire \Q_reg[27]_i_8_n_2 ;
  wire \Q_reg[27]_i_8_n_3 ;
  wire \Q_reg[28]_i_1_n_0 ;
  wire \Q_reg[28]_i_1_n_1 ;
  wire \Q_reg[28]_i_1_n_2 ;
  wire \Q_reg[28]_i_1_n_3 ;
  wire \Q_reg[29]_i_14_n_0 ;
  wire \Q_reg[29]_i_14_n_1 ;
  wire \Q_reg[29]_i_14_n_2 ;
  wire \Q_reg[29]_i_14_n_3 ;
  wire \Q_reg[29]_i_9_n_0 ;
  wire \Q_reg[29]_i_9_n_1 ;
  wire \Q_reg[29]_i_9_n_2 ;
  wire \Q_reg[29]_i_9_n_3 ;
  wire \Q_reg[30]_i_18_n_0 ;
  wire \Q_reg[30]_i_18_n_1 ;
  wire \Q_reg[30]_i_18_n_2 ;
  wire \Q_reg[30]_i_18_n_3 ;
  wire \Q_reg[30]_i_7_n_3 ;
  wire \Q_reg[31]_i_1_n_2 ;
  wire \Q_reg[31]_i_1_n_3 ;
  wire \Q_reg[35]_i_30_n_0 ;
  wire \Q_reg[35]_i_30_n_1 ;
  wire \Q_reg[35]_i_30_n_2 ;
  wire \Q_reg[35]_i_30_n_3 ;
  wire \Q_reg[35]_i_31_n_0 ;
  wire \Q_reg[35]_i_31_n_1 ;
  wire \Q_reg[35]_i_31_n_2 ;
  wire \Q_reg[35]_i_31_n_3 ;
  wire \Q_reg[35]_i_33_n_0 ;
  wire \Q_reg[35]_i_33_n_1 ;
  wire \Q_reg[35]_i_33_n_2 ;
  wire \Q_reg[35]_i_33_n_3 ;
  wire \Q_reg[35]_i_34_n_0 ;
  wire \Q_reg[35]_i_34_n_1 ;
  wire \Q_reg[35]_i_34_n_2 ;
  wire \Q_reg[35]_i_34_n_3 ;
  wire \Q_reg[49]_i_17_n_0 ;
  wire \Q_reg[49]_i_17_n_1 ;
  wire \Q_reg[49]_i_17_n_2 ;
  wire \Q_reg[49]_i_17_n_3 ;
  wire \Q_reg[49]_i_17_n_4 ;
  wire \Q_reg[49]_i_17_n_5 ;
  wire \Q_reg[49]_i_17_n_6 ;
  wire \Q_reg[49]_i_17_n_7 ;
  wire \Q_reg[49]_i_18_n_0 ;
  wire \Q_reg[49]_i_18_n_1 ;
  wire \Q_reg[49]_i_18_n_2 ;
  wire \Q_reg[49]_i_18_n_3 ;
  wire \Q_reg[49]_i_18_n_4 ;
  wire \Q_reg[49]_i_18_n_5 ;
  wire \Q_reg[49]_i_18_n_6 ;
  wire \Q_reg[49]_i_18_n_7 ;
  wire \Q_reg[49]_i_21_n_0 ;
  wire \Q_reg[49]_i_21_n_1 ;
  wire \Q_reg[49]_i_21_n_2 ;
  wire \Q_reg[49]_i_21_n_3 ;
  wire \Q_reg[49]_i_21_n_4 ;
  wire \Q_reg[49]_i_21_n_5 ;
  wire \Q_reg[49]_i_21_n_6 ;
  wire \Q_reg[49]_i_21_n_7 ;
  wire \Q_reg[49]_i_32_n_0 ;
  wire \Q_reg[49]_i_32_n_1 ;
  wire \Q_reg[49]_i_32_n_2 ;
  wire \Q_reg[49]_i_32_n_3 ;
  wire \Q_reg[49]_i_32_n_4 ;
  wire \Q_reg[49]_i_32_n_5 ;
  wire \Q_reg[49]_i_32_n_6 ;
  wire \Q_reg[49]_i_32_n_7 ;
  wire \Q_reg[49]_i_35_n_0 ;
  wire \Q_reg[49]_i_35_n_1 ;
  wire \Q_reg[49]_i_35_n_2 ;
  wire \Q_reg[49]_i_35_n_3 ;
  wire \Q_reg[49]_i_35_n_4 ;
  wire \Q_reg[49]_i_35_n_5 ;
  wire \Q_reg[49]_i_35_n_6 ;
  wire \Q_reg[49]_i_35_n_7 ;
  wire \Q_reg[49]_i_6_n_0 ;
  wire \Q_reg[49]_i_6_n_1 ;
  wire \Q_reg[49]_i_6_n_2 ;
  wire \Q_reg[49]_i_6_n_3 ;
  wire \Q_reg[4]_i_1_n_0 ;
  wire \Q_reg[4]_i_1_n_1 ;
  wire \Q_reg[4]_i_1_n_2 ;
  wire \Q_reg[4]_i_1_n_3 ;
  wire \Q_reg[4]_i_2__0_n_0 ;
  wire \Q_reg[4]_i_2__0_n_1 ;
  wire \Q_reg[4]_i_2__0_n_2 ;
  wire \Q_reg[4]_i_2__0_n_3 ;
  wire \Q_reg[4]_i_2_n_0 ;
  wire \Q_reg[4]_i_2_n_1 ;
  wire \Q_reg[4]_i_2_n_2 ;
  wire \Q_reg[4]_i_2_n_3 ;
  wire \Q_reg[65]_i_6_n_0 ;
  wire \Q_reg[65]_i_6_n_1 ;
  wire \Q_reg[65]_i_6_n_2 ;
  wire \Q_reg[65]_i_6_n_3 ;
  wire \Q_reg[67]_i_2_n_0 ;
  wire \Q_reg[67]_i_2_n_1 ;
  wire \Q_reg[67]_i_2_n_2 ;
  wire \Q_reg[67]_i_2_n_3 ;
  wire \Q_reg[67]_i_3_n_0 ;
  wire \Q_reg[67]_i_3_n_1 ;
  wire \Q_reg[67]_i_3_n_2 ;
  wire \Q_reg[67]_i_3_n_3 ;
  wire \Q_reg[71]_i_2_n_0 ;
  wire \Q_reg[71]_i_2_n_1 ;
  wire \Q_reg[71]_i_2_n_2 ;
  wire \Q_reg[71]_i_2_n_3 ;
  wire \Q_reg[71]_i_3_n_0 ;
  wire \Q_reg[71]_i_3_n_1 ;
  wire \Q_reg[71]_i_3_n_2 ;
  wire \Q_reg[71]_i_3_n_3 ;
  wire \Q_reg[75]_i_2_n_0 ;
  wire \Q_reg[75]_i_2_n_1 ;
  wire \Q_reg[75]_i_2_n_2 ;
  wire \Q_reg[75]_i_2_n_3 ;
  wire \Q_reg[75]_i_3_n_0 ;
  wire \Q_reg[75]_i_3_n_1 ;
  wire \Q_reg[75]_i_3_n_2 ;
  wire \Q_reg[75]_i_3_n_3 ;
  wire \Q_reg[79]_i_2_n_0 ;
  wire \Q_reg[79]_i_2_n_1 ;
  wire \Q_reg[79]_i_2_n_2 ;
  wire \Q_reg[79]_i_2_n_3 ;
  wire \Q_reg[79]_i_3_n_0 ;
  wire \Q_reg[79]_i_3_n_1 ;
  wire \Q_reg[79]_i_3_n_2 ;
  wire \Q_reg[79]_i_3_n_3 ;
  wire \Q_reg[83]_i_2_n_0 ;
  wire \Q_reg[83]_i_2_n_1 ;
  wire \Q_reg[83]_i_2_n_2 ;
  wire \Q_reg[83]_i_2_n_3 ;
  wire \Q_reg[83]_i_3_n_0 ;
  wire \Q_reg[83]_i_3_n_1 ;
  wire \Q_reg[83]_i_3_n_2 ;
  wire \Q_reg[83]_i_3_n_3 ;
  wire \Q_reg[87]_i_2_n_0 ;
  wire \Q_reg[87]_i_2_n_1 ;
  wire \Q_reg[87]_i_2_n_2 ;
  wire \Q_reg[87]_i_2_n_3 ;
  wire \Q_reg[87]_i_3_n_1 ;
  wire \Q_reg[87]_i_3_n_2 ;
  wire \Q_reg[87]_i_3_n_3 ;
  wire \Q_reg[8]_i_1_n_0 ;
  wire \Q_reg[8]_i_1_n_1 ;
  wire \Q_reg[8]_i_1_n_2 ;
  wire \Q_reg[8]_i_1_n_3 ;
  wire \Q_reg[8]_i_2__0_n_0 ;
  wire \Q_reg[8]_i_2__0_n_1 ;
  wire \Q_reg[8]_i_2__0_n_2 ;
  wire \Q_reg[8]_i_2__0_n_3 ;
  wire \Q_reg[8]_i_2_n_0 ;
  wire \Q_reg[8]_i_2_n_1 ;
  wire \Q_reg[8]_i_2_n_2 ;
  wire \Q_reg[8]_i_2_n_3 ;
  wire \Q_reg[9]_i_5_n_1 ;
  wire \Q_reg[9]_i_5_n_2 ;
  wire \Q_reg[9]_i_5_n_3 ;
  wire [4:0]RF_RA1;
  wire [4:0]RF_RA2;
  wire [31:0]RF_RD1;
  wire [31:0]RF_RD1_IBUF;
  wire [31:0]RF_RD2;
  wire [31:0]RF_RD2_IBUF;
  wire [4:0]RF_WA;
  wire [31:0]RF_WD;
  wire RF_WE;
  wire RF_WE_OBUF;
  wire RST0;
  wire RST02_out;
  wire RSTn;
  wire RSTn_IBUF;
  wire [9:0]STALL_COUNTER_D;
  wire STALL_COUNTER_D1;
  wire [9:0]STALL_COUNTER_Q;
  wire STALL_EN;
  wire VCC_2;
  wire WB_CUSTOM_RD;
  wire [31:1]\alu/data0 ;
  wire [31:0]\alu/data1 ;
  wire [31:0]\alu/data2 ;
  wire \alu/data5 ;
  wire \branch_comp/EQ ;
  wire \branch_comp/LT20_in ;
  wire [31:0]\custom_alu/FADD_Q ;
  wire [63:0]\custom_alu/MULT ;
  wire [31:0]\custom_alu/Q ;
  wire [23:1]\custom_alu/fp2int/INT0 ;
  wire \custom_alu/fp2int/INT0_carry__0_n_0 ;
  wire \custom_alu/fp2int/INT0_carry__0_n_1 ;
  wire \custom_alu/fp2int/INT0_carry__0_n_2 ;
  wire \custom_alu/fp2int/INT0_carry__0_n_3 ;
  wire \custom_alu/fp2int/INT0_carry__1_n_0 ;
  wire \custom_alu/fp2int/INT0_carry__1_n_1 ;
  wire \custom_alu/fp2int/INT0_carry__1_n_2 ;
  wire \custom_alu/fp2int/INT0_carry__1_n_3 ;
  wire \custom_alu/fp2int/INT0_carry__2_n_0 ;
  wire \custom_alu/fp2int/INT0_carry__2_n_1 ;
  wire \custom_alu/fp2int/INT0_carry__2_n_2 ;
  wire \custom_alu/fp2int/INT0_carry__2_n_3 ;
  wire \custom_alu/fp2int/INT0_carry__3_n_0 ;
  wire \custom_alu/fp2int/INT0_carry__3_n_1 ;
  wire \custom_alu/fp2int/INT0_carry__3_n_2 ;
  wire \custom_alu/fp2int/INT0_carry__3_n_3 ;
  wire \custom_alu/fp2int/INT0_carry__4_n_0 ;
  wire \custom_alu/fp2int/INT0_carry__4_n_2 ;
  wire \custom_alu/fp2int/INT0_carry__4_n_3 ;
  wire \custom_alu/fp2int/INT0_carry_n_0 ;
  wire \custom_alu/fp2int/INT0_carry_n_1 ;
  wire \custom_alu/fp2int/INT0_carry_n_2 ;
  wire \custom_alu/fp2int/INT0_carry_n_3 ;
  wire [23:0]\custom_alu/fp2int/p_0_in ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[0] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[10] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[11] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[12] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[13] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[14] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[15] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[16] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[17] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[18] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[19] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[1] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[20] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[21] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[22] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[23] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[24] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[25] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[26] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[27] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[28] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[29] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[2] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[30] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[31] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[3] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[4] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[5] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[6] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[7] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[8] ;
  wire \custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[9] ;
  wire [22:1]\custom_alu/fp32_add/data23 ;
  wire [7:0]\custom_alu/fp32_add/exp_a ;
  wire [7:0]\custom_alu/fp32_add/exp_b_add_sub ;
  wire \custom_alu/fp32_add/exp_b_add_sub_carry__0_n_1 ;
  wire \custom_alu/fp32_add/exp_b_add_sub_carry__0_n_2 ;
  wire \custom_alu/fp32_add/exp_b_add_sub_carry__0_n_3 ;
  wire \custom_alu/fp32_add/exp_b_add_sub_carry_n_0 ;
  wire \custom_alu/fp32_add/exp_b_add_sub_carry_n_1 ;
  wire \custom_alu/fp32_add/exp_b_add_sub_carry_n_2 ;
  wire \custom_alu/fp32_add/exp_b_add_sub_carry_n_3 ;
  wire \custom_alu/fp32_add/exp_diff_carry__0_n_1 ;
  wire \custom_alu/fp32_add/exp_diff_carry__0_n_2 ;
  wire \custom_alu/fp32_add/exp_diff_carry__0_n_3 ;
  wire \custom_alu/fp32_add/exp_diff_carry_n_0 ;
  wire \custom_alu/fp32_add/exp_diff_carry_n_1 ;
  wire \custom_alu/fp32_add/exp_diff_carry_n_2 ;
  wire \custom_alu/fp32_add/exp_diff_carry_n_3 ;
  wire [7:0]\custom_alu/fp32_add/exp_sub ;
  wire \custom_alu/fp32_add/op_a2 ;
  wire \custom_alu/fp32_add/op_a2_carry__0_n_0 ;
  wire \custom_alu/fp32_add/op_a2_carry__0_n_1 ;
  wire \custom_alu/fp32_add/op_a2_carry__0_n_2 ;
  wire \custom_alu/fp32_add/op_a2_carry__0_n_3 ;
  wire \custom_alu/fp32_add/op_a2_carry__1_n_0 ;
  wire \custom_alu/fp32_add/op_a2_carry__1_n_1 ;
  wire \custom_alu/fp32_add/op_a2_carry__1_n_2 ;
  wire \custom_alu/fp32_add/op_a2_carry__1_n_3 ;
  wire \custom_alu/fp32_add/op_a2_carry__2_n_1 ;
  wire \custom_alu/fp32_add/op_a2_carry__2_n_2 ;
  wire \custom_alu/fp32_add/op_a2_carry__2_n_3 ;
  wire \custom_alu/fp32_add/op_a2_carry_n_0 ;
  wire \custom_alu/fp32_add/op_a2_carry_n_1 ;
  wire \custom_alu/fp32_add/op_a2_carry_n_2 ;
  wire \custom_alu/fp32_add/op_a2_carry_n_3 ;
  wire [7:0]\custom_alu/fp32_add/p_0_in ;
  wire [6:0]\custom_alu/fp32_add/p_0_in2_in ;
  wire \custom_alu/fp32_add/p_1_in ;
  wire [7:0]\custom_alu/fp32_add/p_1_in__0 ;
  wire [88:1]\custom_alu/fp32_add/p_1_out ;
  wire \custom_alu/fp32_add/pe/exp_sub_carry__0_n_1 ;
  wire \custom_alu/fp32_add/pe/exp_sub_carry__0_n_2 ;
  wire \custom_alu/fp32_add/pe/exp_sub_carry__0_n_3 ;
  wire \custom_alu/fp32_add/pe/exp_sub_carry_n_0 ;
  wire \custom_alu/fp32_add/pe/exp_sub_carry_n_1 ;
  wire \custom_alu/fp32_add/pe/exp_sub_carry_n_2 ;
  wire \custom_alu/fp32_add/pe/exp_sub_carry_n_3 ;
  wire [24:0]\custom_alu/fp32_add/sel0 ;
  wire [24:0]\custom_alu/fp32_add/significand_add0 ;
  wire [23:0]\custom_alu/fp32_add/significand_b_add_sub ;
  wire [24:0]\custom_alu/fp32_add/significand_sub0 ;
  wire [23:0]\custom_alu/fp32_add/significand_sub_complement ;
  wire \custom_alu/fp32_add/significand_sub_complement1 ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[23] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[24] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[25] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[26] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[27] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[28] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[29] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[30] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[31] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[55] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[56] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[57] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[58] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[59] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[60] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[61] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[62] ;
  wire \custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[63] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[23] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[24] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[25] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[26] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[27] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[28] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[29] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[30] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[31] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[55] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[56] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[57] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[58] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[59] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[60] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[61] ;
  wire \custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[62] ;
  wire [24:0]\custom_alu/fp32_mult/PSUM1_2 ;
  wire [31:31]\custom_alu/fp32_mult/a_Q ;
  wire \custom_alu/fp32_mult/exponent_carry__0_n_0 ;
  wire \custom_alu/fp32_mult/exponent_carry__0_n_1 ;
  wire \custom_alu/fp32_mult/exponent_carry__0_n_2 ;
  wire \custom_alu/fp32_mult/exponent_carry__0_n_3 ;
  wire \custom_alu/fp32_mult/exponent_carry__0_n_5 ;
  wire \custom_alu/fp32_mult/exponent_carry__0_n_6 ;
  wire \custom_alu/fp32_mult/exponent_carry__0_n_7 ;
  wire \custom_alu/fp32_mult/exponent_carry__1_n_7 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_0 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_1 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_2 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_3 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_4 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_5 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_6 ;
  wire \custom_alu/fp32_mult/exponent_carry_n_7 ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[0] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[10] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[11] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[12] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[13] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[14] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[15] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[16] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[17] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[18] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[19] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[1] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[20] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[21] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[22] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[23] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[24] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[2] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[3] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[4] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[5] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[6] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[7] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[8] ;
  wire \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[9] ;
  wire [23:0]\custom_alu/fp32_mult/mult24_0/PSUM0__0 ;
  wire [23:0]\custom_alu/fp32_mult/mult24_0/PSUM1__0 ;
  wire [23:0]\custom_alu/fp32_mult/mult24_0/PSUM3__0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[11]_i_2_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[11]_i_3_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[11]_i_4_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[11]_i_5_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[15]_i_2_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[15]_i_3_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[15]_i_4_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[15]_i_5_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[19]_i_2_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[19]_i_3_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[19]_i_4_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[19]_i_5_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[23]_i_2_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[23]_i_3_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[23]_i_4_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[23]_i_5_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[3]_i_2_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[3]_i_3_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[3]_i_4_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[3]_i_5_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[7]_i_2_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[7]_i_3_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[7]_i_4_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q[7]_i_5_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_1 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_2 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_3 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_1 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_2 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_3 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_1 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_2 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_3 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_1 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_2 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_3 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_1 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_2 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_3 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_0 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_1 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_2 ;
  wire \custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_3 ;
  wire \custom_alu/fp32_mult/normalised ;
  wire \custom_alu/fp32_mult/op_a1 ;
  wire \custom_alu/fp32_mult/op_b1 ;
  wire [23:0]\custom_alu/fp32_mult/p_0_in ;
  wire \custom_alu/fp32_mult/p_0_in1_in ;
  wire [47:0]\custom_alu/fp32_mult/p_1_in ;
  wire [22:0]\custom_alu/fp32_mult/product_mantissa ;
  wire [30:1]\custom_alu/int2fp/INT_VAL0 ;
  wire [22:0]\custom_alu/int2fp/INT_VAL1 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[0]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[100]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[101]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[102]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[1]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[2]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[3]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[4]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[5]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[6]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[96]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[97]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[98]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg[99]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__0_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__10_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__11_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__12_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__1_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__2_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__3_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__4_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__5_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__6_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__7_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__8_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate__9_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_gate_n_0 ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[103] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[104] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[105] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[106] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[107] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[108] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[109] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[110] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[111] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[112] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[113] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[114] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[115] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[116] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[117] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[118] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[119] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[120] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[121] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[122] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[123] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[124] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[125] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[126] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[127] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[17] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[18] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[19] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[20] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[21] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[22] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[23] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[49] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[50] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[51] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[52] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[53] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[54] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[55] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[56] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[57] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[58] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[59] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[60] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[61] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[62] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[63] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[64] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[65] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[66] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[67] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[68] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[69] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[70] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[71] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[72] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[73] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[74] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[75] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[76] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[77] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[78] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[79] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[80] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[81] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[82] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[83] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[84] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[85] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[86] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[87] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[88] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[89] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[90] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[91] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[92] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[93] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[94] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[95] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[17] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[18] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[19] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[20] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[21] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[22] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[23] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[49] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[50] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[51] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[52] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[53] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[54] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[55] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[56] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[57] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[58] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[59] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[60] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[61] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[62] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[63] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[64] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[65] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[66] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[67] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[68] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[69] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[70] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[71] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[72] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[73] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[74] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[75] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[76] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[77] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[78] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[79] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[80] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[81] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[82] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[83] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[84] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[85] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[86] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[87] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[88] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[89] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[90] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[91] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[92] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[93] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[94] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[95] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[96] ;
  wire \custom_alu/mult/FF_MULT_1/Q_reg_n_0_[9] ;
  wire [15:0]\custom_alu/mult/PSUM0 ;
  wire [31:7]\custom_alu/mult/PSUM0_1_2_3 ;
  wire [15:0]\custom_alu/mult/PSUM1 ;
  wire [16:0]\custom_alu/mult/PSUM1_2 ;
  wire [15:0]\custom_alu/mult/PSUM2 ;
  wire [15:0]\custom_alu/mult/PSUM3 ;
  wire \custom_alu/mult/Q[11]_i_12_n_0 ;
  wire \custom_alu/mult/Q[11]_i_13_n_0 ;
  wire \custom_alu/mult/Q[11]_i_14_n_0 ;
  wire \custom_alu/mult/Q[11]_i_15_n_0 ;
  wire \custom_alu/mult/Q[11]_i_2_n_0 ;
  wire \custom_alu/mult/Q[11]_i_3_n_0 ;
  wire \custom_alu/mult/Q[11]_i_4_n_0 ;
  wire \custom_alu/mult/Q[11]_i_5_n_0 ;
  wire \custom_alu/mult/Q[15]_i_10_n_0 ;
  wire \custom_alu/mult/Q[15]_i_11_n_0 ;
  wire \custom_alu/mult/Q[15]_i_2_n_0 ;
  wire \custom_alu/mult/Q[15]_i_3_n_0 ;
  wire \custom_alu/mult/Q[15]_i_4_n_0 ;
  wire \custom_alu/mult/Q[15]_i_5_n_0 ;
  wire \custom_alu/mult/Q[15]_i_8_n_0 ;
  wire \custom_alu/mult/Q[15]_i_9_n_0 ;
  wire \custom_alu/mult/Q[19]_i_10_n_0 ;
  wire \custom_alu/mult/Q[19]_i_11_n_0 ;
  wire \custom_alu/mult/Q[19]_i_2_n_0 ;
  wire \custom_alu/mult/Q[19]_i_3_n_0 ;
  wire \custom_alu/mult/Q[19]_i_4_n_0 ;
  wire \custom_alu/mult/Q[19]_i_5_n_0 ;
  wire \custom_alu/mult/Q[19]_i_8_n_0 ;
  wire \custom_alu/mult/Q[19]_i_9_n_0 ;
  wire \custom_alu/mult/Q[23]_i_10_n_0 ;
  wire \custom_alu/mult/Q[23]_i_11_n_0 ;
  wire \custom_alu/mult/Q[23]_i_12_n_0 ;
  wire \custom_alu/mult/Q[23]_i_2_n_0 ;
  wire \custom_alu/mult/Q[23]_i_3_n_0 ;
  wire \custom_alu/mult/Q[23]_i_4_n_0 ;
  wire \custom_alu/mult/Q[23]_i_5_n_0 ;
  wire \custom_alu/mult/Q[23]_i_8_n_0 ;
  wire \custom_alu/mult/Q[23]_i_9_n_0 ;
  wire \custom_alu/mult/Q[27]_i_10_n_0 ;
  wire \custom_alu/mult/Q[27]_i_11_n_0 ;
  wire \custom_alu/mult/Q[27]_i_12_n_0 ;
  wire \custom_alu/mult/Q[27]_i_2_n_0 ;
  wire \custom_alu/mult/Q[27]_i_3_n_0 ;
  wire \custom_alu/mult/Q[27]_i_4_n_0 ;
  wire \custom_alu/mult/Q[27]_i_5_n_0 ;
  wire \custom_alu/mult/Q[27]_i_9_n_0 ;
  wire \custom_alu/mult/Q[31]_i_15_n_0 ;
  wire \custom_alu/mult/Q[31]_i_16_n_0 ;
  wire \custom_alu/mult/Q[31]_i_17_n_0 ;
  wire \custom_alu/mult/Q[31]_i_18_n_0 ;
  wire \custom_alu/mult/Q[31]_i_2_n_0 ;
  wire \custom_alu/mult/Q[31]_i_3_n_0 ;
  wire \custom_alu/mult/Q[31]_i_4_n_0 ;
  wire \custom_alu/mult/Q[31]_i_5_n_0 ;
  wire \custom_alu/mult/Q[35]_i_12_n_0 ;
  wire \custom_alu/mult/Q[35]_i_13_n_0 ;
  wire \custom_alu/mult/Q[35]_i_14_n_0 ;
  wire \custom_alu/mult/Q[35]_i_15_n_0 ;
  wire \custom_alu/mult/Q[3]_i_2_n_0 ;
  wire \custom_alu/mult/Q[3]_i_3_n_0 ;
  wire \custom_alu/mult/Q[3]_i_4_n_0 ;
  wire \custom_alu/mult/Q[3]_i_5_n_0 ;
  wire \custom_alu/mult/Q[5]_i_6_n_0 ;
  wire \custom_alu/mult/Q[5]_i_7_n_0 ;
  wire \custom_alu/mult/Q[5]_i_8_n_0 ;
  wire \custom_alu/mult/Q[5]_i_9_n_0 ;
  wire \custom_alu/mult/Q[7]_i_2_n_0 ;
  wire \custom_alu/mult/Q[7]_i_3_n_0 ;
  wire \custom_alu/mult/Q[7]_i_4_n_0 ;
  wire \custom_alu/mult/Q[7]_i_5_n_0 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[11]_i_1_n_7 ;
  wire \custom_alu/mult/Q_reg[11]_i_8_n_0 ;
  wire \custom_alu/mult/Q_reg[11]_i_8_n_1 ;
  wire \custom_alu/mult/Q_reg[11]_i_8_n_2 ;
  wire \custom_alu/mult/Q_reg[11]_i_8_n_3 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[15]_i_1_n_7 ;
  wire \custom_alu/mult/Q_reg[15]_i_5_n_0 ;
  wire \custom_alu/mult/Q_reg[15]_i_5_n_1 ;
  wire \custom_alu/mult/Q_reg[15]_i_5_n_2 ;
  wire \custom_alu/mult/Q_reg[15]_i_5_n_3 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[19]_i_1_n_7 ;
  wire \custom_alu/mult/Q_reg[19]_i_6_n_0 ;
  wire \custom_alu/mult/Q_reg[19]_i_6_n_1 ;
  wire \custom_alu/mult/Q_reg[19]_i_6_n_2 ;
  wire \custom_alu/mult/Q_reg[19]_i_6_n_3 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[23]_i_1_n_7 ;
  wire \custom_alu/mult/Q_reg[23]_i_4_n_0 ;
  wire \custom_alu/mult/Q_reg[23]_i_4_n_1 ;
  wire \custom_alu/mult/Q_reg[23]_i_4_n_2 ;
  wire \custom_alu/mult/Q_reg[23]_i_4_n_3 ;
  wire \custom_alu/mult/Q_reg[23]_i_5_n_0 ;
  wire \custom_alu/mult/Q_reg[23]_i_5_n_1 ;
  wire \custom_alu/mult/Q_reg[23]_i_5_n_2 ;
  wire \custom_alu/mult/Q_reg[23]_i_5_n_3 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[27]_i_1_n_7 ;
  wire \custom_alu/mult/Q_reg[27]_i_4_n_0 ;
  wire \custom_alu/mult/Q_reg[27]_i_4_n_1 ;
  wire \custom_alu/mult/Q_reg[27]_i_4_n_2 ;
  wire \custom_alu/mult/Q_reg[27]_i_4_n_3 ;
  wire \custom_alu/mult/Q_reg[27]_i_5_n_0 ;
  wire \custom_alu/mult/Q_reg[27]_i_5_n_1 ;
  wire \custom_alu/mult/Q_reg[27]_i_5_n_2 ;
  wire \custom_alu/mult/Q_reg[27]_i_5_n_3 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[31]_i_1_n_7 ;
  wire \custom_alu/mult/Q_reg[31]_i_8_n_0 ;
  wire \custom_alu/mult/Q_reg[31]_i_8_n_1 ;
  wire \custom_alu/mult/Q_reg[31]_i_8_n_2 ;
  wire \custom_alu/mult/Q_reg[31]_i_8_n_3 ;
  wire \custom_alu/mult/Q_reg[31]_i_9_n_0 ;
  wire \custom_alu/mult/Q_reg[31]_i_9_n_1 ;
  wire \custom_alu/mult/Q_reg[31]_i_9_n_2 ;
  wire \custom_alu/mult/Q_reg[31]_i_9_n_3 ;
  wire \custom_alu/mult/Q_reg[32]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[35]_i_5_n_0 ;
  wire \custom_alu/mult/Q_reg[35]_i_5_n_1 ;
  wire \custom_alu/mult/Q_reg[35]_i_5_n_2 ;
  wire \custom_alu/mult/Q_reg[35]_i_5_n_3 ;
  wire \custom_alu/mult/Q_reg[35]_i_6_n_0 ;
  wire \custom_alu/mult/Q_reg[35]_i_6_n_1 ;
  wire \custom_alu/mult/Q_reg[35]_i_6_n_2 ;
  wire \custom_alu/mult/Q_reg[35]_i_6_n_3 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[3]_i_1_n_7 ;
  wire \custom_alu/mult/Q_reg[5]_i_4_n_0 ;
  wire \custom_alu/mult/Q_reg[5]_i_4_n_1 ;
  wire \custom_alu/mult/Q_reg[5]_i_4_n_2 ;
  wire \custom_alu/mult/Q_reg[5]_i_4_n_3 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_0 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_1 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_2 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_3 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_4 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_5 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_6 ;
  wire \custom_alu/mult/Q_reg[7]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[55] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[56] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[57] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[58] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[59] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[60] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[61] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[62] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[63] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM0__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM0__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM1__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM1__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM2__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM2__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_0/PSUM3__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_0/PSUM3__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_0/Q[106]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[106]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[106]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[110]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[110]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[110]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[110]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[114]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[114]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[114]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[114]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[118]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[118]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[118]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[118]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[11]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[11]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[11]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[11]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[122]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[122]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[15]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[15]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[15]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[15]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[3]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[3]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[3]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[3]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[7]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[7]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[7]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_0/Q[7]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[17] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[18] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[19] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[20] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[21] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[22] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[23] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[49] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[50] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[51] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[52] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[53] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[54] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[55] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[56] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[57] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[58] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[59] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[60] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[61] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[62] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[63] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[17] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[18] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[19] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[20] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[21] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[22] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[23] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM0__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM1__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM2__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_1/PSUM3__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_1/Q[11]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[11]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[11]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[11]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[15]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[15]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[15]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[15]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[3]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[3]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[3]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[3]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[74]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[74]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[74]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[78]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[78]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[78]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[78]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[7]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[7]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[7]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[7]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[82]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[82]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[82]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[82]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[86]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[86]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[86]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[86]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[90]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_1/Q[90]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[16]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_1/Q_reg[95]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[17] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[18] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[19] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[20] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[21] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[22] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[23] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[49] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[50] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[51] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[52] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[53] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[54] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[55] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[56] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[57] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[58] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[59] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[60] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[61] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[62] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[63] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[17] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[18] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[19] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[20] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[21] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[22] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[23] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM0__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM1__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM2__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_2/PSUM3__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_2/Q[11]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[11]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[11]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[11]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[15]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[15]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[15]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[15]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[3]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[3]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[3]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[3]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[42]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[42]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[42]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[46]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[46]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[46]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[46]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[50]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[50]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[50]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[50]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[54]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[54]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[54]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[54]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[58]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[58]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[7]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[7]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[7]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_2/Q[7]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[16]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[63]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[17] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[18] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[19] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[20] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[21] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[22] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[23] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[55] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[56] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[57] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[58] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[59] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[60] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[61] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[62] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[63] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[0] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[10] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[11] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[12] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[13] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[14] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[15] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[16] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[1] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[24] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[25] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[26] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[27] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[28] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[29] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[2] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[30] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[31] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[32] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[33] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[34] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[35] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[36] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[37] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[38] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[39] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[3] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[40] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[41] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[42] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[43] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[44] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[45] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[46] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[47] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[48] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[4] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[5] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[6] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[7] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[8] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[9] ;
  wire \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_r_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM0__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM1__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM2__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__0_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__30_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry__2_n_7 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_0 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_1 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_2 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_3 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_4 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_5 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_6 ;
  wire \custom_alu/mult/mult16_3/PSUM3__60_carry_n_7 ;
  wire \custom_alu/mult/mult16_3/Q[10]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[10]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[10]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[11]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[11]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[11]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[11]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[14]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[14]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[14]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[14]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[15]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[15]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[15]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[15]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[18]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[18]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[18]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[18]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[22]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[22]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[22]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[22]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[26]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[26]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[3]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[3]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[3]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[3]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[7]_i_2_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[7]_i_3_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[7]_i_4_n_0 ;
  wire \custom_alu/mult/mult16_3/Q[7]_i_5_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[16]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[31]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_7 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_0 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_1 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_2 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_3 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_4 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_5 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_6 ;
  wire \custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_7 ;
  wire [15:0]\custom_alu/mult/p_0_in ;
  wire [15:0]\custom_alu/mult/p_1_in ;
  wire [31:0]data0;
  wire [31:0]data1;
  wire exp_b_add_sub_carry__0_i_4_n_0;
  wire exp_b_add_sub_carry__0_i_5_n_0;
  wire exp_b_add_sub_carry__0_i_6_n_0;
  wire exp_b_add_sub_carry__0_i_7_n_0;
  wire exp_b_add_sub_carry_i_5_n_0;
  wire exp_b_add_sub_carry_i_6_n_0;
  wire exp_b_add_sub_carry_i_7_n_0;
  wire exp_b_add_sub_carry_i_8_n_0;
  wire exp_diff_carry__0_i_1_n_0;
  wire exp_diff_carry__0_i_2_n_0;
  wire exp_diff_carry__0_i_3_n_0;
  wire exp_diff_carry__0_i_4_n_0;
  wire exp_diff_carry__0_i_5_n_0;
  wire exp_diff_carry__0_i_6_n_0;
  wire exp_diff_carry__0_i_7_n_0;
  wire exp_diff_carry_i_1_n_0;
  wire exp_diff_carry_i_2_n_0;
  wire exp_diff_carry_i_3_n_0;
  wire exp_diff_carry_i_4_n_0;
  wire exp_diff_carry_i_5_n_0;
  wire exp_diff_carry_i_6_n_0;
  wire exp_diff_carry_i_7_n_0;
  wire exp_diff_carry_i_8_n_0;
  wire exp_sub_carry__0_i_1_n_0;
  wire exp_sub_carry__0_i_2_n_0;
  wire exp_sub_carry__0_i_3_n_0;
  wire exp_sub_carry__0_i_4_n_0;
  wire exp_sub_carry__0_i_5_n_0;
  wire exp_sub_carry__0_i_6_n_0;
  wire exp_sub_carry__0_i_7_n_0;
  wire exp_sub_carry__0_i_8_n_0;
  wire exp_sub_carry_i_10_n_0;
  wire exp_sub_carry_i_11_n_0;
  wire exp_sub_carry_i_12_n_0;
  wire exp_sub_carry_i_13_n_0;
  wire exp_sub_carry_i_14_n_0;
  wire exp_sub_carry_i_15_n_0;
  wire exp_sub_carry_i_16_n_0;
  wire exp_sub_carry_i_17_n_0;
  wire exp_sub_carry_i_18_n_0;
  wire exp_sub_carry_i_19_n_0;
  wire exp_sub_carry_i_1_n_0;
  wire exp_sub_carry_i_20_n_0;
  wire exp_sub_carry_i_21_n_0;
  wire exp_sub_carry_i_22_n_0;
  wire exp_sub_carry_i_23_n_0;
  wire exp_sub_carry_i_24_n_0;
  wire exp_sub_carry_i_2_n_0;
  wire exp_sub_carry_i_3_n_0;
  wire exp_sub_carry_i_4_n_0;
  wire exp_sub_carry_i_5_n_0;
  wire exp_sub_carry_i_6_n_0;
  wire exp_sub_carry_i_7_n_0;
  wire exp_sub_carry_i_8_n_0;
  wire exp_sub_carry_i_9_n_0;
  wire exponent_carry__0_i_1_n_0;
  wire exponent_carry__0_i_2_n_0;
  wire exponent_carry__0_i_3_n_0;
  wire exponent_carry__0_i_4_n_0;
  wire exponent_carry__0_i_5_n_0;
  wire exponent_carry__0_i_6_n_0;
  wire exponent_carry__0_i_7_n_0;
  wire exponent_carry__0_i_8_n_0;
  wire exponent_carry__1_i_1_n_0;
  wire exponent_carry_i_10_n_0;
  wire exponent_carry_i_10_n_1;
  wire exponent_carry_i_10_n_2;
  wire exponent_carry_i_10_n_3;
  wire exponent_carry_i_10_n_4;
  wire exponent_carry_i_10_n_5;
  wire exponent_carry_i_10_n_6;
  wire exponent_carry_i_10_n_7;
  wire exponent_carry_i_11_n_0;
  wire exponent_carry_i_11_n_1;
  wire exponent_carry_i_11_n_2;
  wire exponent_carry_i_11_n_3;
  wire exponent_carry_i_11_n_4;
  wire exponent_carry_i_11_n_5;
  wire exponent_carry_i_11_n_6;
  wire exponent_carry_i_11_n_7;
  wire exponent_carry_i_1_n_0;
  wire exponent_carry_i_2_n_0;
  wire exponent_carry_i_3_n_0;
  wire exponent_carry_i_4_n_0;
  wire exponent_carry_i_5_n_0;
  wire exponent_carry_i_6_n_0;
  wire exponent_carry_i_7_n_0;
  wire exponent_carry_i_9_n_0;
  wire exponent_carry_i_9_n_1;
  wire exponent_carry_i_9_n_2;
  wire exponent_carry_i_9_n_3;
  wire exponent_carry_i_9_n_4;
  wire exponent_carry_i_9_n_5;
  wire exponent_carry_i_9_n_6;
  wire exponent_carry_i_9_n_7;
  wire \fp32_add/Q[12]_i_10_n_0 ;
  wire \fp32_add/Q[12]_i_7_n_0 ;
  wire \fp32_add/Q[12]_i_8_n_0 ;
  wire \fp32_add/Q[12]_i_9_n_0 ;
  wire \fp32_add/Q[16]_i_10_n_0 ;
  wire \fp32_add/Q[16]_i_7_n_0 ;
  wire \fp32_add/Q[16]_i_8_n_0 ;
  wire \fp32_add/Q[16]_i_9_n_0 ;
  wire \fp32_add/Q[20]_i_10_n_0 ;
  wire \fp32_add/Q[20]_i_7_n_0 ;
  wire \fp32_add/Q[20]_i_8_n_0 ;
  wire \fp32_add/Q[20]_i_9_n_0 ;
  wire \fp32_add/Q[23]_i_10_n_0 ;
  wire \fp32_add/Q[23]_i_8_n_0 ;
  wire \fp32_add/Q[23]_i_9_n_0 ;
  wire \fp32_add/Q[4]_i_10_n_0 ;
  wire \fp32_add/Q[4]_i_7_n_0 ;
  wire \fp32_add/Q[4]_i_8_n_0 ;
  wire \fp32_add/Q[4]_i_9_n_0 ;
  wire \fp32_add/Q[67]_i_4_n_0 ;
  wire \fp32_add/Q[67]_i_5_n_0 ;
  wire \fp32_add/Q[67]_i_6_n_0 ;
  wire \fp32_add/Q[67]_i_7_n_0 ;
  wire \fp32_add/Q[71]_i_4_n_0 ;
  wire \fp32_add/Q[71]_i_5_n_0 ;
  wire \fp32_add/Q[71]_i_6_n_0 ;
  wire \fp32_add/Q[71]_i_7_n_0 ;
  wire \fp32_add/Q[75]_i_4_n_0 ;
  wire \fp32_add/Q[75]_i_5_n_0 ;
  wire \fp32_add/Q[75]_i_6_n_0 ;
  wire \fp32_add/Q[75]_i_7_n_0 ;
  wire \fp32_add/Q[79]_i_4_n_0 ;
  wire \fp32_add/Q[79]_i_5_n_0 ;
  wire \fp32_add/Q[79]_i_6_n_0 ;
  wire \fp32_add/Q[79]_i_7_n_0 ;
  wire \fp32_add/Q[83]_i_4_n_0 ;
  wire \fp32_add/Q[83]_i_5_n_0 ;
  wire \fp32_add/Q[83]_i_6_n_0 ;
  wire \fp32_add/Q[83]_i_7_n_0 ;
  wire \fp32_add/Q[87]_i_5_n_0 ;
  wire \fp32_add/Q[87]_i_6_n_0 ;
  wire \fp32_add/Q[87]_i_7_n_0 ;
  wire \fp32_add/Q[8]_i_10_n_0 ;
  wire \fp32_add/Q[8]_i_7_n_0 ;
  wire \fp32_add/Q[8]_i_8_n_0 ;
  wire \fp32_add/Q[8]_i_9_n_0 ;
  wire \fp32_mult/mult24_0/Q[16]_i_14_n_0 ;
  wire \fp32_mult/mult24_0/Q[16]_i_15_n_0 ;
  wire \fp32_mult/mult24_0/Q[16]_i_16_n_0 ;
  wire \fp32_mult/mult24_0/Q[16]_i_17_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_24_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_25_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_26_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_27_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_28_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_29_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_30_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_31_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_37_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_38_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_39_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_40_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_41_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_42_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_43_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_44_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_45_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_46_n_0 ;
  wire \fp32_mult/mult24_0/Q[49]_i_47_n_0 ;
  wire \fp32_mult/mult24_0/exponent_carry_i_12_n_0 ;
  wire \fp32_mult/mult24_0/exponent_carry_i_13_n_0 ;
  wire op_a2_carry__0_i_1_n_0;
  wire op_a2_carry__0_i_2_n_0;
  wire op_a2_carry__0_i_3_n_0;
  wire op_a2_carry__0_i_4_n_0;
  wire op_a2_carry__0_i_5_n_0;
  wire op_a2_carry__0_i_6_n_0;
  wire op_a2_carry__0_i_7_n_0;
  wire op_a2_carry__0_i_8_n_0;
  wire op_a2_carry__1_i_1_n_0;
  wire op_a2_carry__1_i_2_n_0;
  wire op_a2_carry__1_i_3_n_0;
  wire op_a2_carry__1_i_4_n_0;
  wire op_a2_carry__1_i_5_n_0;
  wire op_a2_carry__1_i_6_n_0;
  wire op_a2_carry__1_i_7_n_0;
  wire op_a2_carry__1_i_8_n_0;
  wire op_a2_carry__2_i_1_n_0;
  wire op_a2_carry__2_i_2_n_0;
  wire op_a2_carry__2_i_3_n_0;
  wire op_a2_carry__2_i_4_n_0;
  wire op_a2_carry__2_i_5_n_0;
  wire op_a2_carry__2_i_6_n_0;
  wire op_a2_carry__2_i_7_n_0;
  wire op_a2_carry__2_i_8_n_0;
  wire op_a2_carry_i_1_n_0;
  wire op_a2_carry_i_2_n_0;
  wire op_a2_carry_i_3_n_0;
  wire op_a2_carry_i_4_n_0;
  wire op_a2_carry_i_5_n_0;
  wire op_a2_carry_i_6_n_0;
  wire op_a2_carry_i_7_n_0;
  wire op_a2_carry_i_8_n_0;
  wire op_a2_carry_i_9_n_0;
  wire [0:0]p_0_in;
  wire \stall_generator/CUSTOM_STALL ;
  wire \stall_generator/LU_HAZARD1 ;
  wire \stall_generator/LU_HAZARD17_out ;
  wire [3:0]\NLW_custom_alu/fp2int/INT0_carry__4_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM0__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM0__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM1__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM1__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM2__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM2__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM3__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_0/PSUM3__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM0__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM0__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM1__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM1__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM2__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM2__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM3__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_1/PSUM3__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM0__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM0__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM1__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM1__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM2__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM2__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM3__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_2/PSUM3__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM0__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM0__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM1__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM1__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM2__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM2__30_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM3__0_carry__1_CO_UNCONNECTED ;
  wire [3:0]\NLW_custom_alu/mult/mult16_3/PSUM3__30_carry__1_CO_UNCONNECTED ;

  BUFG CLK_IBUF_BUFG_inst
       (.I(CLK_IBUF),
        .O(CLK_IBUF_BUFG));
  IBUF CLK_IBUF_inst
       (.I(CLK),
        .O(CLK_IBUF));
  OBUF \CRF_RA1_OBUF[0]_inst 
       (.I(CRF_RA1_OBUF[0]),
        .O(CRF_RA1[0]));
  OBUF \CRF_RA1_OBUF[1]_inst 
       (.I(CRF_RA1_OBUF[1]),
        .O(CRF_RA1[1]));
  OBUF \CRF_RA1_OBUF[2]_inst 
       (.I(CRF_RA1_OBUF[2]),
        .O(CRF_RA1[2]));
  OBUF \CRF_RA1_OBUF[3]_inst 
       (.I(CRF_RA1_OBUF[3]),
        .O(CRF_RA1[3]));
  OBUF \CRF_RA1_OBUF[4]_inst 
       (.I(CRF_RA1_OBUF[4]),
        .O(CRF_RA1[4]));
  OBUF \CRF_RA2_OBUF[0]_inst 
       (.I(CRF_RA2_OBUF[0]),
        .O(CRF_RA2[0]));
  OBUF \CRF_RA2_OBUF[1]_inst 
       (.I(CRF_RA2_OBUF[1]),
        .O(CRF_RA2[1]));
  OBUF \CRF_RA2_OBUF[2]_inst 
       (.I(CRF_RA2_OBUF[2]),
        .O(CRF_RA2[2]));
  OBUF \CRF_RA2_OBUF[3]_inst 
       (.I(CRF_RA2_OBUF[3]),
        .O(CRF_RA2[3]));
  OBUF \CRF_RA2_OBUF[4]_inst 
       (.I(CRF_RA2_OBUF[4]),
        .O(CRF_RA2[4]));
  IBUF \CRF_RD1_IBUF[0]_inst 
       (.I(CRF_RD1[0]),
        .O(CRF_RD1_IBUF[0]));
  IBUF \CRF_RD1_IBUF[10]_inst 
       (.I(CRF_RD1[10]),
        .O(CRF_RD1_IBUF[10]));
  IBUF \CRF_RD1_IBUF[11]_inst 
       (.I(CRF_RD1[11]),
        .O(CRF_RD1_IBUF[11]));
  IBUF \CRF_RD1_IBUF[12]_inst 
       (.I(CRF_RD1[12]),
        .O(CRF_RD1_IBUF[12]));
  IBUF \CRF_RD1_IBUF[13]_inst 
       (.I(CRF_RD1[13]),
        .O(CRF_RD1_IBUF[13]));
  IBUF \CRF_RD1_IBUF[14]_inst 
       (.I(CRF_RD1[14]),
        .O(CRF_RD1_IBUF[14]));
  IBUF \CRF_RD1_IBUF[15]_inst 
       (.I(CRF_RD1[15]),
        .O(CRF_RD1_IBUF[15]));
  IBUF \CRF_RD1_IBUF[16]_inst 
       (.I(CRF_RD1[16]),
        .O(CRF_RD1_IBUF[16]));
  IBUF \CRF_RD1_IBUF[17]_inst 
       (.I(CRF_RD1[17]),
        .O(CRF_RD1_IBUF[17]));
  IBUF \CRF_RD1_IBUF[18]_inst 
       (.I(CRF_RD1[18]),
        .O(CRF_RD1_IBUF[18]));
  IBUF \CRF_RD1_IBUF[19]_inst 
       (.I(CRF_RD1[19]),
        .O(CRF_RD1_IBUF[19]));
  IBUF \CRF_RD1_IBUF[1]_inst 
       (.I(CRF_RD1[1]),
        .O(CRF_RD1_IBUF[1]));
  IBUF \CRF_RD1_IBUF[20]_inst 
       (.I(CRF_RD1[20]),
        .O(CRF_RD1_IBUF[20]));
  IBUF \CRF_RD1_IBUF[21]_inst 
       (.I(CRF_RD1[21]),
        .O(CRF_RD1_IBUF[21]));
  IBUF \CRF_RD1_IBUF[22]_inst 
       (.I(CRF_RD1[22]),
        .O(CRF_RD1_IBUF[22]));
  IBUF \CRF_RD1_IBUF[23]_inst 
       (.I(CRF_RD1[23]),
        .O(CRF_RD1_IBUF[23]));
  IBUF \CRF_RD1_IBUF[24]_inst 
       (.I(CRF_RD1[24]),
        .O(CRF_RD1_IBUF[24]));
  IBUF \CRF_RD1_IBUF[25]_inst 
       (.I(CRF_RD1[25]),
        .O(CRF_RD1_IBUF[25]));
  IBUF \CRF_RD1_IBUF[26]_inst 
       (.I(CRF_RD1[26]),
        .O(CRF_RD1_IBUF[26]));
  IBUF \CRF_RD1_IBUF[27]_inst 
       (.I(CRF_RD1[27]),
        .O(CRF_RD1_IBUF[27]));
  IBUF \CRF_RD1_IBUF[28]_inst 
       (.I(CRF_RD1[28]),
        .O(CRF_RD1_IBUF[28]));
  IBUF \CRF_RD1_IBUF[29]_inst 
       (.I(CRF_RD1[29]),
        .O(CRF_RD1_IBUF[29]));
  IBUF \CRF_RD1_IBUF[2]_inst 
       (.I(CRF_RD1[2]),
        .O(CRF_RD1_IBUF[2]));
  IBUF \CRF_RD1_IBUF[30]_inst 
       (.I(CRF_RD1[30]),
        .O(CRF_RD1_IBUF[30]));
  IBUF \CRF_RD1_IBUF[31]_inst 
       (.I(CRF_RD1[31]),
        .O(CRF_RD1_IBUF[31]));
  IBUF \CRF_RD1_IBUF[3]_inst 
       (.I(CRF_RD1[3]),
        .O(CRF_RD1_IBUF[3]));
  IBUF \CRF_RD1_IBUF[4]_inst 
       (.I(CRF_RD1[4]),
        .O(CRF_RD1_IBUF[4]));
  IBUF \CRF_RD1_IBUF[5]_inst 
       (.I(CRF_RD1[5]),
        .O(CRF_RD1_IBUF[5]));
  IBUF \CRF_RD1_IBUF[6]_inst 
       (.I(CRF_RD1[6]),
        .O(CRF_RD1_IBUF[6]));
  IBUF \CRF_RD1_IBUF[7]_inst 
       (.I(CRF_RD1[7]),
        .O(CRF_RD1_IBUF[7]));
  IBUF \CRF_RD1_IBUF[8]_inst 
       (.I(CRF_RD1[8]),
        .O(CRF_RD1_IBUF[8]));
  IBUF \CRF_RD1_IBUF[9]_inst 
       (.I(CRF_RD1[9]),
        .O(CRF_RD1_IBUF[9]));
  IBUF \CRF_RD2_IBUF[0]_inst 
       (.I(CRF_RD2[0]),
        .O(CRF_RD2_IBUF[0]));
  IBUF \CRF_RD2_IBUF[10]_inst 
       (.I(CRF_RD2[10]),
        .O(CRF_RD2_IBUF[10]));
  IBUF \CRF_RD2_IBUF[11]_inst 
       (.I(CRF_RD2[11]),
        .O(CRF_RD2_IBUF[11]));
  IBUF \CRF_RD2_IBUF[12]_inst 
       (.I(CRF_RD2[12]),
        .O(CRF_RD2_IBUF[12]));
  IBUF \CRF_RD2_IBUF[13]_inst 
       (.I(CRF_RD2[13]),
        .O(CRF_RD2_IBUF[13]));
  IBUF \CRF_RD2_IBUF[14]_inst 
       (.I(CRF_RD2[14]),
        .O(CRF_RD2_IBUF[14]));
  IBUF \CRF_RD2_IBUF[15]_inst 
       (.I(CRF_RD2[15]),
        .O(CRF_RD2_IBUF[15]));
  IBUF \CRF_RD2_IBUF[16]_inst 
       (.I(CRF_RD2[16]),
        .O(CRF_RD2_IBUF[16]));
  IBUF \CRF_RD2_IBUF[17]_inst 
       (.I(CRF_RD2[17]),
        .O(CRF_RD2_IBUF[17]));
  IBUF \CRF_RD2_IBUF[18]_inst 
       (.I(CRF_RD2[18]),
        .O(CRF_RD2_IBUF[18]));
  IBUF \CRF_RD2_IBUF[19]_inst 
       (.I(CRF_RD2[19]),
        .O(CRF_RD2_IBUF[19]));
  IBUF \CRF_RD2_IBUF[1]_inst 
       (.I(CRF_RD2[1]),
        .O(CRF_RD2_IBUF[1]));
  IBUF \CRF_RD2_IBUF[20]_inst 
       (.I(CRF_RD2[20]),
        .O(CRF_RD2_IBUF[20]));
  IBUF \CRF_RD2_IBUF[21]_inst 
       (.I(CRF_RD2[21]),
        .O(CRF_RD2_IBUF[21]));
  IBUF \CRF_RD2_IBUF[22]_inst 
       (.I(CRF_RD2[22]),
        .O(CRF_RD2_IBUF[22]));
  IBUF \CRF_RD2_IBUF[23]_inst 
       (.I(CRF_RD2[23]),
        .O(CRF_RD2_IBUF[23]));
  IBUF \CRF_RD2_IBUF[24]_inst 
       (.I(CRF_RD2[24]),
        .O(CRF_RD2_IBUF[24]));
  IBUF \CRF_RD2_IBUF[25]_inst 
       (.I(CRF_RD2[25]),
        .O(CRF_RD2_IBUF[25]));
  IBUF \CRF_RD2_IBUF[26]_inst 
       (.I(CRF_RD2[26]),
        .O(CRF_RD2_IBUF[26]));
  IBUF \CRF_RD2_IBUF[27]_inst 
       (.I(CRF_RD2[27]),
        .O(CRF_RD2_IBUF[27]));
  IBUF \CRF_RD2_IBUF[28]_inst 
       (.I(CRF_RD2[28]),
        .O(CRF_RD2_IBUF[28]));
  IBUF \CRF_RD2_IBUF[29]_inst 
       (.I(CRF_RD2[29]),
        .O(CRF_RD2_IBUF[29]));
  IBUF \CRF_RD2_IBUF[2]_inst 
       (.I(CRF_RD2[2]),
        .O(CRF_RD2_IBUF[2]));
  IBUF \CRF_RD2_IBUF[30]_inst 
       (.I(CRF_RD2[30]),
        .O(CRF_RD2_IBUF[30]));
  IBUF \CRF_RD2_IBUF[31]_inst 
       (.I(CRF_RD2[31]),
        .O(CRF_RD2_IBUF[31]));
  IBUF \CRF_RD2_IBUF[3]_inst 
       (.I(CRF_RD2[3]),
        .O(CRF_RD2_IBUF[3]));
  IBUF \CRF_RD2_IBUF[4]_inst 
       (.I(CRF_RD2[4]),
        .O(CRF_RD2_IBUF[4]));
  IBUF \CRF_RD2_IBUF[5]_inst 
       (.I(CRF_RD2[5]),
        .O(CRF_RD2_IBUF[5]));
  IBUF \CRF_RD2_IBUF[6]_inst 
       (.I(CRF_RD2[6]),
        .O(CRF_RD2_IBUF[6]));
  IBUF \CRF_RD2_IBUF[7]_inst 
       (.I(CRF_RD2[7]),
        .O(CRF_RD2_IBUF[7]));
  IBUF \CRF_RD2_IBUF[8]_inst 
       (.I(CRF_RD2[8]),
        .O(CRF_RD2_IBUF[8]));
  IBUF \CRF_RD2_IBUF[9]_inst 
       (.I(CRF_RD2[9]),
        .O(CRF_RD2_IBUF[9]));
  OBUF \CRF_WA_OBUF[0]_inst 
       (.I(CRF_WA_OBUF[0]),
        .O(CRF_WA[0]));
  OBUF \CRF_WA_OBUF[1]_inst 
       (.I(CRF_WA_OBUF[1]),
        .O(CRF_WA[1]));
  OBUF \CRF_WA_OBUF[2]_inst 
       (.I(CRF_WA_OBUF[2]),
        .O(CRF_WA[2]));
  OBUF \CRF_WA_OBUF[3]_inst 
       (.I(CRF_WA_OBUF[3]),
        .O(CRF_WA[3]));
  OBUF \CRF_WA_OBUF[4]_inst 
       (.I(CRF_WA_OBUF[4]),
        .O(CRF_WA[4]));
  OBUF \CRF_WD_OBUF[0]_inst 
       (.I(CRF_WD_OBUF[0]),
        .O(CRF_WD[0]));
  OBUF \CRF_WD_OBUF[10]_inst 
       (.I(CRF_WD_OBUF[10]),
        .O(CRF_WD[10]));
  OBUF \CRF_WD_OBUF[11]_inst 
       (.I(CRF_WD_OBUF[11]),
        .O(CRF_WD[11]));
  OBUF \CRF_WD_OBUF[12]_inst 
       (.I(CRF_WD_OBUF[12]),
        .O(CRF_WD[12]));
  OBUF \CRF_WD_OBUF[13]_inst 
       (.I(CRF_WD_OBUF[13]),
        .O(CRF_WD[13]));
  OBUF \CRF_WD_OBUF[14]_inst 
       (.I(CRF_WD_OBUF[14]),
        .O(CRF_WD[14]));
  OBUF \CRF_WD_OBUF[15]_inst 
       (.I(CRF_WD_OBUF[15]),
        .O(CRF_WD[15]));
  OBUF \CRF_WD_OBUF[16]_inst 
       (.I(CRF_WD_OBUF[16]),
        .O(CRF_WD[16]));
  OBUF \CRF_WD_OBUF[17]_inst 
       (.I(CRF_WD_OBUF[17]),
        .O(CRF_WD[17]));
  OBUF \CRF_WD_OBUF[18]_inst 
       (.I(CRF_WD_OBUF[18]),
        .O(CRF_WD[18]));
  OBUF \CRF_WD_OBUF[19]_inst 
       (.I(CRF_WD_OBUF[19]),
        .O(CRF_WD[19]));
  OBUF \CRF_WD_OBUF[1]_inst 
       (.I(CRF_WD_OBUF[1]),
        .O(CRF_WD[1]));
  OBUF \CRF_WD_OBUF[20]_inst 
       (.I(CRF_WD_OBUF[20]),
        .O(CRF_WD[20]));
  OBUF \CRF_WD_OBUF[21]_inst 
       (.I(CRF_WD_OBUF[21]),
        .O(CRF_WD[21]));
  OBUF \CRF_WD_OBUF[22]_inst 
       (.I(CRF_WD_OBUF[22]),
        .O(CRF_WD[22]));
  OBUF \CRF_WD_OBUF[23]_inst 
       (.I(CRF_WD_OBUF[23]),
        .O(CRF_WD[23]));
  OBUF \CRF_WD_OBUF[24]_inst 
       (.I(CRF_WD_OBUF[24]),
        .O(CRF_WD[24]));
  OBUF \CRF_WD_OBUF[25]_inst 
       (.I(CRF_WD_OBUF[25]),
        .O(CRF_WD[25]));
  OBUF \CRF_WD_OBUF[26]_inst 
       (.I(CRF_WD_OBUF[26]),
        .O(CRF_WD[26]));
  OBUF \CRF_WD_OBUF[27]_inst 
       (.I(CRF_WD_OBUF[27]),
        .O(CRF_WD[27]));
  OBUF \CRF_WD_OBUF[28]_inst 
       (.I(CRF_WD_OBUF[28]),
        .O(CRF_WD[28]));
  OBUF \CRF_WD_OBUF[29]_inst 
       (.I(CRF_WD_OBUF[29]),
        .O(CRF_WD[29]));
  OBUF \CRF_WD_OBUF[2]_inst 
       (.I(CRF_WD_OBUF[2]),
        .O(CRF_WD[2]));
  OBUF \CRF_WD_OBUF[30]_inst 
       (.I(CRF_WD_OBUF[30]),
        .O(CRF_WD[30]));
  OBUF \CRF_WD_OBUF[31]_inst 
       (.I(CRF_WD_OBUF[31]),
        .O(CRF_WD[31]));
  OBUF \CRF_WD_OBUF[3]_inst 
       (.I(CRF_WD_OBUF[3]),
        .O(CRF_WD[3]));
  OBUF \CRF_WD_OBUF[4]_inst 
       (.I(CRF_WD_OBUF[4]),
        .O(CRF_WD[4]));
  OBUF \CRF_WD_OBUF[5]_inst 
       (.I(CRF_WD_OBUF[5]),
        .O(CRF_WD[5]));
  OBUF \CRF_WD_OBUF[6]_inst 
       (.I(CRF_WD_OBUF[6]),
        .O(CRF_WD[6]));
  OBUF \CRF_WD_OBUF[7]_inst 
       (.I(CRF_WD_OBUF[7]),
        .O(CRF_WD[7]));
  OBUF \CRF_WD_OBUF[8]_inst 
       (.I(CRF_WD_OBUF[8]),
        .O(CRF_WD[8]));
  OBUF \CRF_WD_OBUF[9]_inst 
       (.I(CRF_WD_OBUF[9]),
        .O(CRF_WD[9]));
  OBUF CRF_WE_OBUF_inst
       (.I(CRF_WE_OBUF),
        .O(CRF_WE));
  LUT2 #(
    .INIT(4'h8)) 
    CRF_WE_OBUF_inst_i_1
       (.I0(WB_CUSTOM_RD),
        .I1(MEM_WB_Q),
        .O(CRF_WE_OBUF));
  OBUF \D_MEM_ADDR_OBUF[0]_inst 
       (.I(D_MEM_ADDR_OBUF[0]),
        .O(D_MEM_ADDR[0]));
  LUT6 #(
    .INIT(64'hFFFFABAAAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[0]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[0]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[0]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[0]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[0]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[0]));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_10 
       (.I0(ALU_DIN2[1]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN1[0]),
        .I4(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_19_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_20_n_0 ),
        .I3(ALU_DIN2[2]),
        .I4(\D_MEM_ADDR_OBUF[8]_inst_i_16_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[0]_inst_i_14_n_0 ),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_12 
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN1[8]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[16]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[0]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_12_n_0 ));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \D_MEM_ADDR_OBUF[0]_inst_i_13 
       (.CI(\D_MEM_ADDR_OBUF[0]_inst_i_15_n_0 ),
        .CO({\alu/data5 ,\D_MEM_ADDR_OBUF[0]_inst_i_13_n_1 ,\D_MEM_ADDR_OBUF[0]_inst_i_13_n_2 ,\D_MEM_ADDR_OBUF[0]_inst_i_13_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\D_MEM_ADDR_OBUF[0]_inst_i_16_n_0 ,op_a2_carry__2_i_2_n_0,op_a2_carry__2_i_3_n_0,op_a2_carry__2_i_4_n_0}),
        .S({\D_MEM_ADDR_OBUF[0]_inst_i_17_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_19_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_20_n_0 }));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_14 
       (.I0(ALU_DIN1[16]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[0]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_14_n_0 ));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \D_MEM_ADDR_OBUF[0]_inst_i_15 
       (.CI(\D_MEM_ADDR_OBUF[0]_inst_i_21_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[0]_inst_i_15_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_15_n_1 ,\D_MEM_ADDR_OBUF[0]_inst_i_15_n_2 ,\D_MEM_ADDR_OBUF[0]_inst_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI({op_a2_carry__1_i_1_n_0,op_a2_carry__1_i_2_n_0,op_a2_carry__1_i_3_n_0,op_a2_carry__1_i_4_n_0}),
        .S({\D_MEM_ADDR_OBUF[0]_inst_i_22_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_23_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_24_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_25_n_0 }));
  LUT6 #(
    .INIT(64'h54045404FD5D5404)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_16 
       (.I0(\Q[63]_i_1__1_n_0 ),
        .I1(EX_RF_RD2[31]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(ID_EX_Q[110]),
        .I4(ALU_DIN2[30]),
        .I5(ALU_DIN1[30]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hE21D00000000E21D)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_17 
       (.I0(EX_RF_RD2[31]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[110]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[30]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_18 
       (.I0(ALU_DIN1[29]),
        .I1(ID_EX_Q[108]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[29]),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[28]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_19 
       (.I0(ALU_DIN1[27]),
        .I1(ID_EX_Q[106]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[27]),
        .I4(ALU_DIN1[26]),
        .I5(ALU_DIN2[26]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_2 
       (.I0(ID_EX_Q[126]),
        .I1(ID_EX_Q[125]),
        .I2(\alu/data1 [0]),
        .I3(ID_EX_Q[123]),
        .I4(\alu/data2 [0]),
        .I5(ID_EX_Q[122]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_20 
       (.I0(ALU_DIN1[25]),
        .I1(ID_EX_Q[104]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[25]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[24]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_20_n_0 ));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \D_MEM_ADDR_OBUF[0]_inst_i_21 
       (.CI(\D_MEM_ADDR_OBUF[0]_inst_i_26_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[0]_inst_i_21_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_21_n_1 ,\D_MEM_ADDR_OBUF[0]_inst_i_21_n_2 ,\D_MEM_ADDR_OBUF[0]_inst_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI({op_a2_carry__0_i_1_n_0,op_a2_carry__0_i_2_n_0,op_a2_carry__0_i_3_n_0,op_a2_carry__0_i_4_n_0}),
        .S({\D_MEM_ADDR_OBUF[0]_inst_i_27_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_28_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_29_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_30_n_0 }));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_22 
       (.I0(ALU_DIN1[23]),
        .I1(ID_EX_Q[102]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[23]),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[22]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_23 
       (.I0(ALU_DIN1[21]),
        .I1(ID_EX_Q[100]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[21]),
        .I4(ALU_DIN1[20]),
        .I5(ALU_DIN2[20]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_24 
       (.I0(ALU_DIN1[19]),
        .I1(ID_EX_Q[98]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[19]),
        .I4(ALU_DIN1[18]),
        .I5(ALU_DIN2[18]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_25 
       (.I0(ALU_DIN1[17]),
        .I1(ID_EX_Q[96]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[17]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[16]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_25_n_0 ));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \D_MEM_ADDR_OBUF[0]_inst_i_26 
       (.CI(\<const0> ),
        .CO({\D_MEM_ADDR_OBUF[0]_inst_i_26_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_26_n_1 ,\D_MEM_ADDR_OBUF[0]_inst_i_26_n_2 ,\D_MEM_ADDR_OBUF[0]_inst_i_26_n_3 }),
        .CYINIT(\<const0> ),
        .DI({op_a2_carry_i_1_n_0,op_a2_carry_i_2_n_0,op_a2_carry_i_3_n_0,op_a2_carry_i_4_n_0}),
        .S({\D_MEM_ADDR_OBUF[0]_inst_i_31_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_32_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_33_n_0 ,\D_MEM_ADDR_OBUF[0]_inst_i_34_n_0 }));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_27 
       (.I0(ALU_DIN1[15]),
        .I1(ID_EX_Q[94]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[15]),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[14]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_28 
       (.I0(ALU_DIN1[13]),
        .I1(ID_EX_Q[92]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[13]),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[12]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_29 
       (.I0(ALU_DIN1[11]),
        .I1(ID_EX_Q[90]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[11]),
        .I4(ALU_DIN1[10]),
        .I5(ALU_DIN2[10]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h020202022A002AAA)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(ALU_DIN1[0]),
        .I3(ID_EX_Q[114]),
        .I4(ID_EX_Q[79]),
        .I5(ID_EX_Q[115]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_30 
       (.I0(ALU_DIN1[9]),
        .I1(ID_EX_Q[88]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[9]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[8]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_31 
       (.I0(ALU_DIN1[7]),
        .I1(ID_EX_Q[86]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[7]),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[6]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h9099900009000999)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_32 
       (.I0(ALU_DIN1[5]),
        .I1(ALU_DIN2[5]),
        .I2(ID_EX_Q[130]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[4]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_33 
       (.I0(ID_EX_Q[129]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[3]),
        .I3(ALU_DIN2[3]),
        .I4(ALU_DIN1[2]),
        .I5(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h9099900009000999)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_34 
       (.I0(ALU_DIN2[0]),
        .I1(ALU_DIN1[0]),
        .I2(ID_EX_Q[127]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[1]),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_4 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[0]),
        .I4(ALU_DIN1[0]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAEEAAAA)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[0]_inst_i_7_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[0]_inst_i_8_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[1]_inst_i_10_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_6 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[0]_inst_i_9_n_0 ),
        .I2(ID_EX_Q[121]),
        .I3(\D_MEM_ADDR_OBUF[0]_inst_i_10_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBB888B8)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[1]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[0]_inst_i_11_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[2]_inst_i_10_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[6]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[1]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_16_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[0]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h888EEE8EAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[0]_inst_i_9 
       (.I0(\alu/data5 ),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I4(ID_EX_Q[110]),
        .I5(ID_EX_Q[120]),
        .O(\D_MEM_ADDR_OBUF[0]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[10]_inst 
       (.I(D_MEM_ADDR_OBUF[10]),
        .O(D_MEM_ADDR[10]));
  LUT6 #(
    .INIT(64'hFF10FFFFFF100000)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[10]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[10]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[10]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[10]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[10]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[10]));
  LUT6 #(
    .INIT(64'h4D48FFFF4D480000)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_10 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[18]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[10]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_11 
       (.I0(ALU_DIN1[3]),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[7]),
        .I4(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_12 
       (.I0(ALU_DIN1[26]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[10]),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_2 
       (.I0(ID_EX_Q[89]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[10]),
        .I3(ALU_DIN2[10]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_3 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[10]),
        .I4(ALU_DIN1[10]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4540)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[11]_inst_i_12_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[10]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[10]_inst_i_8_n_0 ),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hB800)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[10]_inst_i_9_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[11]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_6 
       (.I0(\alu/data0 [10]),
        .I1(ID_EX_Q[125]),
        .I2(\alu/data1 [10]),
        .I3(ID_EX_Q[123]),
        .I4(ID_EX_Q[122]),
        .I5(\alu/data2 [10]),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[14]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[10]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_27_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[12]_inst_i_14_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEAEAAAEAEAAAAAAA)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(ID_EX_Q[117]),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[11]_inst_i_11_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[9]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \D_MEM_ADDR_OBUF[10]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[10]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[12]_inst_i_12_n_0 ),
        .I2(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[10]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[11]_inst 
       (.I(D_MEM_ADDR_OBUF[11]),
        .O(D_MEM_ADDR[11]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[11]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[11]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[11]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[11]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[11]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[11]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[11]));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[11]_inst_i_21_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_13_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[11]_inst_i_22_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_13 
       (.I0(ID_EX_Q[137]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[11]),
        .I3(ID_EX_Q[90]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[11]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_14 
       (.I0(ID_EX_Q[136]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[10]),
        .I3(ID_EX_Q[89]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[10]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_15 
       (.I0(ID_EX_Q[135]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[9]),
        .I3(ID_EX_Q[88]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[9]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_16 
       (.I0(ID_EX_Q[134]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[8]),
        .I3(ID_EX_Q[87]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[8]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_17 
       (.I0(EX_RF_RD2[11]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[90]),
        .I3(EX_RF_RD1[11]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[137]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_18 
       (.I0(EX_RF_RD2[10]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[89]),
        .I3(EX_RF_RD1[10]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[136]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_19 
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[88]),
        .I3(EX_RF_RD1[9]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[135]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_2 
       (.I0(\alu/data2 [11]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [11]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [11]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_20 
       (.I0(EX_RF_RD2[8]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[87]),
        .I3(EX_RF_RD1[8]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[134]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_21 
       (.I0(ALU_DIN1[4]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[0]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[8]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_22 
       (.I0(ALU_DIN1[23]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[11]_inst_i_23_n_0 ),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[7]_inst_i_24_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_23 
       (.I0(ID_EX_Q[157]),
        .I1(EX_RF_RD1[31]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ID_EX_Q[141]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I5(EX_RF_RD1[15]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hD100FFFF)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[12]_inst_i_9_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[11]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[12]_inst_i_10_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[11]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[11]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[12]_inst_i_11_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[11]),
        .I4(ALU_DIN1[11]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[11]_inst_i_7 
       (.I0(ID_EX_Q[90]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[11]),
        .I3(ALU_DIN2[11]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[11]_inst_i_7_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[11]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[7]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[11]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[11]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[11]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[11:8]),
        .O(\alu/data2 [11:8]),
        .S({\D_MEM_ADDR_OBUF[11]_inst_i_13_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_14_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_15_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_16_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[11]_inst_i_9 
       (.CI(\D_MEM_ADDR_OBUF[7]_inst_i_9_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[11]_inst_i_9_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_9_n_1 ,\D_MEM_ADDR_OBUF[11]_inst_i_9_n_2 ,\D_MEM_ADDR_OBUF[11]_inst_i_9_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[11:8]),
        .O(\alu/data1 [11:8]),
        .S({\D_MEM_ADDR_OBUF[11]_inst_i_17_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_19_n_0 ,\D_MEM_ADDR_OBUF[11]_inst_i_20_n_0 }));
  OBUF \D_MEM_ADDR_OBUF[12]_inst 
       (.I(D_MEM_ADDR_OBUF[12]),
        .O(D_MEM_ADDR[12]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[12]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[12]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[12]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[12]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[12]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[12]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[12]));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[14]_inst_i_13_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[12]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_25_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[14]_inst_i_12_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_27_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[12]_inst_i_14_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF5F5FFFF303F)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_12 
       (.I0(ALU_DIN1[5]),
        .I1(ALU_DIN1[1]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[9]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_13 
       (.I0(ALU_DIN1[24]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[16]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[8]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4D48FFFF4D480000)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_14 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[20]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[4]_inst_i_19_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_2 
       (.I0(\alu/data2 [12]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [12]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [12]),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h08A8FFFF)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[13]_inst_i_8_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[12]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[13]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[12]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF470047FF)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_11_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[12]_inst_i_11_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN1[12]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_7 
       (.I0(ID_EX_Q[91]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[12]),
        .I3(ALU_DIN2[12]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_7_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[12]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[8]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[12]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[12]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[12]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[12]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/data0 [12:9]),
        .S(ID_EX_Q[138:135]));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[12]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[12]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[14]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[12]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[13]_inst 
       (.I(D_MEM_ADDR_OBUF[13]),
        .O(D_MEM_ADDR[13]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[13]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[13]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[13]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[13]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[13]));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_15_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_29_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_16_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000A0A0000CFC0)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_12 
       (.I0(ALU_DIN1[6]),
        .I1(ALU_DIN1[2]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[10]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_13 
       (.I0(ALU_DIN1[25]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[17]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[9]_inst_i_16_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F00FB0B0F00F808)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_14 
       (.I0(ALU_DIN1[27]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[19]),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h3F00FB0B3F00F808)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_15 
       (.I0(ALU_DIN1[23]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[15]),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4D48FFFF4D480000)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_16 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[21]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[13]_inst_i_17_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_17 
       (.I0(ALU_DIN1[29]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[13]),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_2 
       (.I0(\alu/data2 [13]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [13]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [13]),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h80A2FFFF)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_8_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[14]_inst_i_8_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[14]_inst_i_10_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[13]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FF4747)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_11_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[14]_inst_i_9_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[13]),
        .I4(ALU_DIN1[13]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_7 
       (.I0(ID_EX_Q[92]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[13]),
        .I3(ALU_DIN2[13]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_31_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[13]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_30_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[13]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[13]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[14]_inst 
       (.I(D_MEM_ADDR_OBUF[14]),
        .O(D_MEM_ADDR[14]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[14]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[14]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[14]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[14]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[14]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[14]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[14]));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[16]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[14]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFCC47FF47)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_11 
       (.I0(ALU_DIN1[7]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[11]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[3]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4D48FFFF4D480000)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_12 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[22]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[4]_inst_i_17_n_0 ),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_13 
       (.I0(ALU_DIN1[26]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[18]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[9]_inst_i_14_n_0 ),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_2 
       (.I0(\alu/data2 [14]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [14]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [14]),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[14]_inst_i_8_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_15_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEAFFEAEAAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_14_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_12_n_0 ),
        .I5(ALU_DIN2[0]),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAFBFBFB)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_5 
       (.I0(ALU_DIN2[0]),
        .I1(\D_MEM_ADDR_OBUF[14]_inst_i_9_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[14]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[14]),
        .I4(ALU_DIN1[14]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_7 
       (.I0(ID_EX_Q[93]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[14]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[14]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[16]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[14]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_25_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[14]_inst_i_12_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_26_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_27_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[14]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[15]_inst 
       (.I(D_MEM_ADDR_OBUF[15]),
        .O(D_MEM_ADDR[15]));
  LUT6 #(
    .INIT(64'hFFFFBBBAAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[15]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_24_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_25_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_26_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_27_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_11 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_28_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_29_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[13]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_13 
       (.I0(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I1(ID_EX_Q[117]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_14 
       (.I0(\D_MEM_ADDR_OBUF[17]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_30_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_14_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_15 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_31_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[17]_inst_i_10_n_0 ),
        .I2(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_16 
       (.I0(EX_RF_RD2[15]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[94]),
        .I3(EX_RF_RD1[15]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[141]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_17 
       (.I0(EX_RF_RD2[14]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[93]),
        .I3(EX_RF_RD1[14]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[140]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_18 
       (.I0(EX_RF_RD2[13]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[92]),
        .I3(EX_RF_RD1[13]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[139]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_19 
       (.I0(EX_RF_RD2[12]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[91]),
        .I3(EX_RF_RD1[12]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[138]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_2 
       (.I0(\alu/data0 [15]),
        .I1(ID_EX_Q[125]),
        .I2(\alu/data1 [15]),
        .I3(ID_EX_Q[123]),
        .I4(\alu/data2 [15]),
        .I5(ID_EX_Q[122]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_20 
       (.I0(ID_EX_Q[141]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[15]),
        .I3(ID_EX_Q[94]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[15]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_21 
       (.I0(ID_EX_Q[140]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[14]),
        .I3(ID_EX_Q[93]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[14]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_22 
       (.I0(ID_EX_Q[139]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[13]),
        .I3(ID_EX_Q[92]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[13]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_23 
       (.I0(ID_EX_Q[138]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[12]),
        .I3(ID_EX_Q[91]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[12]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0F00FB0B0F00F808)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_24 
       (.I0(ALU_DIN1[30]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[22]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0F00FB0B0F00F808)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_25 
       (.I0(ALU_DIN1[26]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[18]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0F00FB0B0F00F808)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_26 
       (.I0(ALU_DIN1[28]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[20]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0F00FB0B0F00F808)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_27 
       (.I0(ALU_DIN1[24]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[16]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0F00FB0B0F00F808)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_28 
       (.I0(ALU_DIN1[29]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[21]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0F00FB0B0F00F808)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_29 
       (.I0(ALU_DIN1[25]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[17]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEAAE)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_9_n_0 ),
        .I1(ID_EX_Q[118]),
        .I2(ALU_DIN1[15]),
        .I3(ALU_DIN2[15]),
        .I4(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_30 
       (.I0(ALU_DIN1[27]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[19]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_32_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_31 
       (.I0(ALU_DIN1[0]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[8]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_33_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_31_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_32 
       (.I0(ALU_DIN1[23]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[15]),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2FFE200)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_33 
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[12]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_33_n_0 ));
  LUT4 #(
    .INIT(16'h2320)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_10_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[16]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_14_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h7400)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_6 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_15_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[16]_inst_i_8_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_6_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[15]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[11]_inst_i_9_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[15]_inst_i_7_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[15]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[15]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[15:12]),
        .O(\alu/data1 [15:12]),
        .S({\D_MEM_ADDR_OBUF[15]_inst_i_16_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_17_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_19_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[15]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[11]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[15]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[15]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[15]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[15:12]),
        .O(\alu/data2 [15:12]),
        .S({\D_MEM_ADDR_OBUF[15]_inst_i_20_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_21_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_22_n_0 ,\D_MEM_ADDR_OBUF[15]_inst_i_23_n_0 }));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[15]_inst_i_9 
       (.I0(ID_EX_Q[94]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[15]),
        .I3(ALU_DIN2[15]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[15]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[16]_inst 
       (.I(D_MEM_ADDR_OBUF[16]),
        .O(D_MEM_ADDR[16]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[16]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[16]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[16]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[16]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[16]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[16]));
  LUT6 #(
    .INIT(64'h4040404444444044)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_10 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_10_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[17]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_11 
       (.I0(ALU_DIN1[1]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[9]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[16]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h88888888B8BBB888)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[16]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[24]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[16]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1D001DFF)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_13 
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[13]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBB888B8)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_14 
       (.I0(ALU_DIN1[28]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(EX_RF_RD1[20]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[146]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_2 
       (.I0(\alu/data2 [16]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [16]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [16]),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[16]_inst_i_8_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[17]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFD55555)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[17]_inst_i_8_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[16]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[16]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[16]),
        .I4(ALU_DIN1[16]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_6 
       (.I0(ID_EX_Q[95]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[16]),
        .I3(ALU_DIN2[16]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_6_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[16]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[12]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[16]_inst_i_7_n_0 ,\D_MEM_ADDR_OBUF[16]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[16]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[16]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/data0 [16:13]),
        .S(ID_EX_Q[142:139]));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT3 #(
    .INIT(8'h74)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[16]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[18]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[16]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[18]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[16]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[16]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[17]_inst 
       (.I(D_MEM_ADDR_OBUF[17]),
        .O(D_MEM_ADDR[17]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[17]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[17]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[17]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[17]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[17]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[17]));
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_10 
       (.I0(ALU_DIN1[2]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[10]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[17]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_11 
       (.I0(ALU_DIN1[29]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[21]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[17]_inst_i_14_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_28_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_29_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_26_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[13]_inst_i_14_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1D001DFF)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_13 
       (.I0(EX_RF_RD1[6]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[132]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[14]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2FFE200)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_14 
       (.I0(EX_RF_RD1[25]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[151]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[17]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_2 
       (.I0(\alu/data2 [17]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [17]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [17]),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8A80FFFF)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[17]_inst_i_7_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[18]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5F5D555)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[18]_inst_i_8_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[17]_inst_i_8_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[17]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN1[17]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_6 
       (.I0(ID_EX_Q[96]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[17]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'h74)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[17]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[19]_inst_i_20_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[19]_inst_i_21_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[17]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4044404040444444)) 
    \D_MEM_ADDR_OBUF[17]_inst_i_9 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[18]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[17]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[17]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[18]_inst 
       (.I(D_MEM_ADDR_OBUF[18]),
        .O(D_MEM_ADDR[18]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[18]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[18]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[18]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[18]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[18]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[18]));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_10 
       (.I0(ALU_DIN1[11]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[3]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[18]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_11 
       (.I0(ALU_DIN1[30]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[22]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[18]_inst_i_14_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_28_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_26_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_24_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_25_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2FFE200)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_13 
       (.I0(EX_RF_RD1[7]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[133]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[15]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2FFE200)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_14 
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[18]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_2 
       (.I0(\alu/data2 [18]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [18]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [18]),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8A80FFFF)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[18]_inst_i_7_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[19]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5D555D5)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[18]_inst_i_8_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[19]_inst_i_10_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[18]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[18]),
        .I4(ALU_DIN1[18]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_6 
       (.I0(ID_EX_Q[97]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[18]),
        .I3(ALU_DIN2[18]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[18]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[20]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[20]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[18]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4044404040444444)) 
    \D_MEM_ADDR_OBUF[18]_inst_i_9 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[19]_inst_i_22_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[18]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[18]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[19]_inst 
       (.I(D_MEM_ADDR_OBUF[19]),
        .O(D_MEM_ADDR[19]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[19]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[19]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[19]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[19]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[19]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[19]));
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[21]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[19]_inst_i_21_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4044404040444444)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_11 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[20]_inst_i_13_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[19]_inst_i_22_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_12 
       (.I0(ID_EX_Q[145]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[19]),
        .I3(ID_EX_Q[98]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[19]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_13 
       (.I0(ID_EX_Q[144]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[18]),
        .I3(ID_EX_Q[97]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[18]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_14 
       (.I0(ID_EX_Q[143]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[17]),
        .I3(ID_EX_Q[96]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[17]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_15 
       (.I0(ID_EX_Q[142]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[16]),
        .I3(ID_EX_Q[95]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[16]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_16 
       (.I0(EX_RF_RD2[19]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[98]),
        .I3(EX_RF_RD1[19]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[145]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_17 
       (.I0(EX_RF_RD2[18]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[97]),
        .I3(EX_RF_RD1[18]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[144]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_18 
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[96]),
        .I3(EX_RF_RD1[17]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[143]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_19 
       (.I0(EX_RF_RD2[16]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[95]),
        .I3(EX_RF_RD1[16]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[142]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_2 
       (.I0(\alu/data2 [19]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [19]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [19]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_20 
       (.I0(ALU_DIN1[4]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[12]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[23]_inst_i_29_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h3022FFFF30220000)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_21 
       (.I0(ALU_DIN1[23]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[19]_inst_i_23_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_22 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_24_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_28_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_26_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[13]_inst_i_14_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2FFE200)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_23 
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[19]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hA808FFFF)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[20]_inst_i_8_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[19]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5DD5555)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[19]_inst_i_10_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[20]_inst_i_9_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[19]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[19]),
        .I4(ALU_DIN1[19]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_6 
       (.I0(ID_EX_Q[98]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[19]),
        .I3(ALU_DIN2[19]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_6_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[19]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[15]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[19]_inst_i_7_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[19]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[19]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[19:16]),
        .O(\alu/data2 [19:16]),
        .S({\D_MEM_ADDR_OBUF[19]_inst_i_12_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_13_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_14_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_15_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[19]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[15]_inst_i_7_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[19]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[19]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[19]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[19:16]),
        .O(\alu/data1 [19:16]),
        .S({\D_MEM_ADDR_OBUF[19]_inst_i_16_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_17_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[19]_inst_i_19_n_0 }));
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[19]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[19]_inst_i_20_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[21]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[19]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[1]_inst 
       (.I(D_MEM_ADDR_OBUF[1]),
        .O(D_MEM_ADDR[1]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[1]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[1]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[1]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[1]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[1]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[1]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[1]));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[7]_inst_i_25_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_30_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_15_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[1]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_31_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[1]_inst_i_14_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_12 
       (.I0(ALU_DIN1[26]),
        .I1(ALU_DIN1[10]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[18]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[2]),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_13 
       (.I0(ALU_DIN1[25]),
        .I1(ALU_DIN1[9]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[17]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[1]),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_14 
       (.I0(\D_MEM_ADDR_OBUF[5]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_21_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[1]_inst_i_15_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_15 
       (.I0(ALU_DIN1[17]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[1]),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_2 
       (.I0(\alu/data2 [1]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [1]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [1]),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h04070000FFFFFFFF)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[1]_inst_i_8_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(ALU_DIN2[1]),
        .I3(\D_MEM_ADDR_OBUF[2]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[1]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[1]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[1]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[2]_inst_i_7_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN1[1]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_7 
       (.I0(ID_EX_Q[80]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[1]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFABFB)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_8 
       (.I0(ALU_DIN2[2]),
        .I1(EX_RF_RD1[0]),
        .I2(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I3(ID_EX_Q[126]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[1]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[6]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[1]_inst_i_12_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[8]_inst_i_14_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_16_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[1]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[20]_inst 
       (.I(D_MEM_ADDR_OBUF[20]),
        .O(D_MEM_ADDR[20]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[20]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[20]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[20]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[20]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[20]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[20]));
  LUT6 #(
    .INIT(64'h4044404040444444)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_10 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[21]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[20]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_11 
       (.I0(ALU_DIN1[5]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[13]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[24]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_12 
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[28]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[20]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_13 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_17_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_24_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_28_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_26_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_2 
       (.I0(\alu/data2 [20]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [20]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [20]),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8A80FFFF)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[20]_inst_i_8_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[21]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5D555D5)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[20]_inst_i_9_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[21]_inst_i_8_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[20]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN1[20]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_6 
       (.I0(ID_EX_Q[99]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[20]),
        .I3(ALU_DIN2[20]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_6_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[20]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[16]_inst_i_7_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[20]_inst_i_7_n_0 ,\D_MEM_ADDR_OBUF[20]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[20]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[20]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/data0 [20:17]),
        .S(ID_EX_Q[146:143]));
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[20]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[22]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[20]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[22]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[20]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[20]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[21]_inst 
       (.I(D_MEM_ADDR_OBUF[21]),
        .O(D_MEM_ADDR[21]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[21]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[21]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[21]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[21]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[21]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[21]));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_10 
       (.I0(ALU_DIN1[6]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[14]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[25]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_11 
       (.I0(ALU_DIN1[25]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[29]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[21]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_24_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[15]_inst_i_28_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_25_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[23]_inst_i_26_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_2 
       (.I0(\alu/data2 [21]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [21]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [21]),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA808FFFF)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[22]_inst_i_7_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[21]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5F5D555)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[22]_inst_i_8_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[21]_inst_i_8_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[21]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[21]),
        .I4(ALU_DIN1[21]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_6 
       (.I0(ID_EX_Q[100]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[21]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[21]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[23]_inst_i_22_n_0 ),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_23_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[21]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4040404444444044)) 
    \D_MEM_ADDR_OBUF[21]_inst_i_9 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[21]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[22]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[21]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[22]_inst 
       (.I(D_MEM_ADDR_OBUF[22]),
        .O(D_MEM_ADDR[22]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[22]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[22]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[22]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[22]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[22]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[22]));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_10 
       (.I0(ALU_DIN1[7]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[15]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[26]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_11 
       (.I0(ALU_DIN1[26]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[30]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[22]),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_27_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[23]_inst_i_28_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_17_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[15]_inst_i_24_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_2 
       (.I0(\alu/data2 [22]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [22]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [22]),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8A80FFFF)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[22]_inst_i_7_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5D555D5)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[22]_inst_i_8_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[23]_inst_i_10_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[22]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[22]),
        .I4(ALU_DIN1[22]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_6 
       (.I0(ID_EX_Q[101]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[22]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[24]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[28]_inst_i_11_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[22]_inst_i_10_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[24]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[22]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4040404444444044)) 
    \D_MEM_ADDR_OBUF[22]_inst_i_9 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[22]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[23]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[22]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[23]_inst 
       (.I(D_MEM_ADDR_OBUF[23]),
        .O(D_MEM_ADDR[23]));
  LUT6 #(
    .INIT(64'h88888888AAAA88A8)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[23]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[23]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_5_n_0 ),
        .I4(ID_EX_Q[118]),
        .I5(\D_MEM_ADDR_OBUF[23]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[23]));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[25]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[23]_inst_i_23_n_0 ),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_16_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[23]_inst_i_24_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_25_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[23]_inst_i_26_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_16_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_17_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_27_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[23]_inst_i_28_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_13 
       (.I0(ID_EX_Q[102]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN2[23]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_14 
       (.I0(ID_EX_Q[149]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[23]),
        .I3(ID_EX_Q[102]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[23]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_15 
       (.I0(ID_EX_Q[148]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[22]),
        .I3(ID_EX_Q[101]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[22]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_16 
       (.I0(ID_EX_Q[147]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[21]),
        .I3(ID_EX_Q[100]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[21]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_17 
       (.I0(ID_EX_Q[146]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[20]),
        .I3(ID_EX_Q[99]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[20]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_18 
       (.I0(EX_RF_RD2[23]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[102]),
        .I3(EX_RF_RD1[23]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[149]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_19 
       (.I0(EX_RF_RD2[22]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[101]),
        .I3(EX_RF_RD1[22]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[148]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_2 
       (.I0(\alu/data2 [23]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [23]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [23]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_20 
       (.I0(EX_RF_RD2[21]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[100]),
        .I3(EX_RF_RD1[21]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[147]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_21 
       (.I0(EX_RF_RD2[20]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[99]),
        .I3(EX_RF_RD1[20]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[146]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h88B8BBBB88B88888)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_22 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_29_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[12]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[27]_inst_i_23_n_0 ),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0033000000B800B8)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_23 
       (.I0(ALU_DIN1[27]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[23]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h10F110E0)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_24 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[25]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h10F110E0)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_25 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[27]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h00F0F0E2)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_26 
       (.I0(ALU_DIN1[23]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[5]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h10F110E0)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_27 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[28]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h10F110E0)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_28 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[24]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_29 
       (.I0(ALU_DIN1[8]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[0]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[16]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h8A80FFFF)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[23]_inst_i_9_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[24]_inst_i_8_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[24]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_10_n_0 ),
        .I4(ID_EX_Q[117]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4040404444444044)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_5 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_11_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[23]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEAAE)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_6 
       (.I0(\D_MEM_ADDR_OBUF[23]_inst_i_13_n_0 ),
        .I1(ID_EX_Q[118]),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN2[23]),
        .I4(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_6_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[23]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[19]_inst_i_7_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[23]_inst_i_7_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[23]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[23]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[23:20]),
        .O(\alu/data2 [23:20]),
        .S({\D_MEM_ADDR_OBUF[23]_inst_i_14_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_15_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_16_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_17_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[23]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[19]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[23]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[23]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[23]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[23:20]),
        .O(\alu/data1 [23:20]),
        .S({\D_MEM_ADDR_OBUF[23]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_19_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_20_n_0 ,\D_MEM_ADDR_OBUF[23]_inst_i_21_n_0 }));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[23]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[25]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[29]_inst_i_14_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_22_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[23]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[24]_inst 
       (.I(D_MEM_ADDR_OBUF[24]),
        .O(D_MEM_ADDR[24]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[24]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[24]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[24]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[24]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[24]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[24]));
  LUT6 #(
    .INIT(64'h4040404444444044)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_10 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[23]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[25]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_11 
       (.I0(ALU_DIN1[9]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[1]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[17]),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00000B08)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_12 
       (.I0(ALU_DIN1[28]),
        .I1(ALU_DIN2[2]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN1[24]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_2 
       (.I0(\alu/data2 [24]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [24]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [24]),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[24]_inst_i_8_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[25]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5DD5555)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[24]_inst_i_9_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[25]_inst_i_8_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[24]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[24]),
        .I4(ALU_DIN1[24]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_6 
       (.I0(ID_EX_Q[103]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[24]),
        .I3(ALU_DIN2[24]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_6_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[24]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[20]_inst_i_7_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[24]_inst_i_7_n_0 ,\D_MEM_ADDR_OBUF[24]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[24]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[24]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/data0 [24:21]),
        .S(ID_EX_Q[150:147]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[24]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[28]_inst_i_11_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_13_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_20_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[24]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[24]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[24]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[25]_inst 
       (.I(D_MEM_ADDR_OBUF[25]),
        .O(D_MEM_ADDR[25]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[25]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[25]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[25]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[25]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[25]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[25]));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_10 
       (.I0(ALU_DIN1[10]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[2]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[18]),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00000B08)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_11 
       (.I0(ALU_DIN1[29]),
        .I1(ALU_DIN2[2]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN1[25]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_16_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[23]_inst_i_24_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_20_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_2 
       (.I0(\alu/data2 [25]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [25]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [25]),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[25]_inst_i_7_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5DD5555)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[25]_inst_i_8_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_8_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[25]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN1[25]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_6 
       (.I0(ID_EX_Q[104]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[25]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[25]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[29]_inst_i_14_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[27]_inst_i_21_n_0 ),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[27]_inst_i_22_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[25]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4044404040444444)) 
    \D_MEM_ADDR_OBUF[25]_inst_i_9 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_10_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[25]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[25]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[26]_inst 
       (.I(D_MEM_ADDR_OBUF[26]),
        .O(D_MEM_ADDR[26]));
  LUT6 #(
    .INIT(64'h88888888AAAA88A8)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[26]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_5_n_0 ),
        .I4(ID_EX_Q[118]),
        .I5(\D_MEM_ADDR_OBUF[26]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[26]));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_16_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_17_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_18_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_19_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_20_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_12 
       (.I0(ID_EX_Q[105]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[26]),
        .I3(ALU_DIN2[26]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_13 
       (.I0(ALU_DIN1[11]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[3]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[19]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00000B08)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_14 
       (.I0(ALU_DIN1[30]),
        .I1(ALU_DIN2[2]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN1[26]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_15 
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN2[24]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN2[29]),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_27_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h10F110E0)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_16 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[30]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h10F110E0)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_17 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[26]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0100FF010100FE00)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_18 
       (.I0(ALU_DIN2[2]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[28]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0100FF010100FE00)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_19 
       (.I0(ALU_DIN2[2]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[29]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_2 
       (.I0(\alu/data2 [26]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [26]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [26]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0300FF010300FE00)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_20 
       (.I0(ALU_DIN2[2]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[27]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_7_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[27]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[27]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_8_n_0 ),
        .I4(ID_EX_Q[117]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4040404444444044)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_5 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_10_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[26]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEAAE)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_6 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_12_n_0 ),
        .I1(ID_EX_Q[118]),
        .I2(ALU_DIN1[26]),
        .I3(ALU_DIN2[26]),
        .I4(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_30_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[26]_inst_i_13_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_20_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(ALU_DIN1[28]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN2[2]),
        .I4(ALU_DIN2[1]),
        .I5(\D_MEM_ADDR_OBUF[26]_inst_i_14_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \D_MEM_ADDR_OBUF[26]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_15_n_0 ),
        .I1(ALU_DIN2[27]),
        .I2(ALU_DIN2[19]),
        .I3(ALU_DIN2[14]),
        .I4(ALU_DIN2[8]),
        .I5(\D_MEM_ADDR_OBUF[31]_inst_i_29_n_0 ),
        .O(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[27]_inst 
       (.I(D_MEM_ADDR_OBUF[27]),
        .O(D_MEM_ADDR[27]));
  LUT6 #(
    .INIT(64'h888888888888AAA8)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[27]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[27]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[27]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[118]),
        .I4(\D_MEM_ADDR_OBUF[27]_inst_i_5_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[27]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[27]));
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(ALU_DIN1[29]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN2[2]),
        .I4(ALU_DIN2[1]),
        .I5(\D_MEM_ADDR_OBUF[27]_inst_i_22_n_0 ),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_11 
       (.I0(ALU_DIN1[30]),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[28]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4044404040444444)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_12 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[28]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[26]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_13 
       (.I0(ID_EX_Q[153]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[27]),
        .I3(ID_EX_Q[106]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[27]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_14 
       (.I0(ID_EX_Q[152]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[26]),
        .I3(ID_EX_Q[105]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[26]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_15 
       (.I0(ID_EX_Q[151]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[25]),
        .I3(ID_EX_Q[104]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[25]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_16 
       (.I0(ID_EX_Q[150]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[24]),
        .I3(ID_EX_Q[103]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[24]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_17 
       (.I0(EX_RF_RD2[27]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[106]),
        .I3(EX_RF_RD1[27]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[153]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_18 
       (.I0(EX_RF_RD2[26]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[105]),
        .I3(EX_RF_RD1[26]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[152]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_19 
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[104]),
        .I3(EX_RF_RD1[25]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[151]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_2 
       (.I0(\alu/data2 [27]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [27]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [27]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_20 
       (.I0(EX_RF_RD2[24]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[103]),
        .I3(EX_RF_RD1[24]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[150]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_21 
       (.I0(ALU_DIN1[12]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[27]_inst_i_23_n_0 ),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[31]_inst_i_22_n_0 ),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h00000B08)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_22 
       (.I0(PSUM3__0_carry__0_i_10__2_n_0),
        .I1(ALU_DIN2[2]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN1[27]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_23 
       (.I0(ID_EX_Q[130]),
        .I1(EX_RF_RD1[4]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ID_EX_Q[146]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I5(EX_RF_RD1[20]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[27]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[28]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5DD5555)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_4 
       (.I0(ID_EX_Q[117]),
        .I1(\D_MEM_ADDR_OBUF[27]_inst_i_10_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[27]_inst_i_11_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[27]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_5 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[27]),
        .I4(ALU_DIN1[27]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_6 
       (.I0(ID_EX_Q[106]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[27]),
        .I3(ALU_DIN2[27]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_6_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[27]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[23]_inst_i_7_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[27]_inst_i_7_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[27]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[27]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[27:24]),
        .O(\alu/data2 [27:24]),
        .S({\D_MEM_ADDR_OBUF[27]_inst_i_13_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_14_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_15_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_16_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[27]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[23]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[27]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[27]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[27]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ALU_DIN1[27:24]),
        .O(\alu/data1 [27:24]),
        .S({\D_MEM_ADDR_OBUF[27]_inst_i_17_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_19_n_0 ,\D_MEM_ADDR_OBUF[27]_inst_i_20_n_0 }));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[27]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_24_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[27]_inst_i_21_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[27]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[28]_inst 
       (.I(D_MEM_ADDR_OBUF[28]),
        .O(D_MEM_ADDR[28]));
  LUT5 #(
    .INIT(32'h8888888A)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[28]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[28]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[28]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[28]));
  LUT6 #(
    .INIT(64'hAEAEAEAAAAAAAEAA)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_10 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[28]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_11 
       (.I0(ALU_DIN1[13]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[5]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[21]),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[30]_inst_i_15_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[26]_inst_i_18_n_0 ),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_2 
       (.I0(\alu/data2 [28]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [28]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [28]),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA280FFFF)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[28]_inst_i_7_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[29]_inst_i_8_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h90FF000090FF90FF)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_4 
       (.I0(ALU_DIN1[28]),
        .I1(ALU_DIN2[28]),
        .I2(ID_EX_Q[118]),
        .I3(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[28]_inst_i_9_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[28]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_5 
       (.I0(ID_EX_Q[107]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[28]),
        .I3(ALU_DIN2[28]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_5_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[28]_inst_i_6 
       (.CI(\D_MEM_ADDR_OBUF[24]_inst_i_7_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[28]_inst_i_6_n_0 ,\D_MEM_ADDR_OBUF[28]_inst_i_6_n_1 ,\D_MEM_ADDR_OBUF[28]_inst_i_6_n_2 ,\D_MEM_ADDR_OBUF[28]_inst_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/data0 [28:25]),
        .S(ID_EX_Q[154:151]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_30_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[30]_inst_i_20_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_33_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_8 
       (.I0(ID_EX_Q[118]),
        .I1(ID_EX_Q[117]),
        .I2(ID_EX_Q[116]),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hEAEFFFFFAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[28]_inst_i_9 
       (.I0(ID_EX_Q[118]),
        .I1(\D_MEM_ADDR_OBUF[29]_inst_i_17_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[27]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I5(ID_EX_Q[117]),
        .O(\D_MEM_ADDR_OBUF[28]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[29]_inst 
       (.I(D_MEM_ADDR_OBUF[29]),
        .O(D_MEM_ADDR[29]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[29]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[29]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[29]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[29]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[29]));
  LUT6 #(
    .INIT(64'h02A2FFFF02A20000)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_10 
       (.I0(\Q[63]_i_1__1_n_0 ),
        .I1(EX_RF_RD2[5]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(ID_EX_Q[84]),
        .I4(ALU_DIN2[1]),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_15_n_0 ),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I1(ID_EX_Q[116]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFEEFFFFAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_12 
       (.I0(ID_EX_Q[118]),
        .I1(\D_MEM_ADDR_OBUF[29]_inst_i_17_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_11_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I5(ID_EX_Q[117]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_13 
       (.I0(ID_EX_Q[117]),
        .I1(ID_EX_Q[116]),
        .I2(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_14 
       (.I0(ALU_DIN1[14]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[6]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[22]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h03F3000057F70000)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_15 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(EX_RF_RD2[5]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(ID_EX_Q[84]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h10F110E0)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_16 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[29]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F7)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_17 
       (.I0(\Q[63]_i_1__1_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[29]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_2 
       (.I0(\alu/data2 [29]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [29]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [29]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA808FFFF)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[30]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[29]_inst_i_8_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00E2)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_9_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[29]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[29]_inst_i_11_n_0 ),
        .I4(ID_EX_Q[117]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0EFE)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_5 
       (.I0(ID_EX_Q[116]),
        .I1(ID_EX_Q[117]),
        .I2(ID_EX_Q[118]),
        .I3(ALU_DIN2[29]),
        .I4(ALU_DIN1[29]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_6 
       (.I0(ID_EX_Q[108]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[29]),
        .I3(ALU_DIN2[29]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_7 
       (.I0(ID_EX_Q[121]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[119]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_24_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_22_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_23_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00F0BBBB00F08888)) 
    \D_MEM_ADDR_OBUF[29]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[29]_inst_i_15_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN2[2]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_16_n_0 ),
        .O(\D_MEM_ADDR_OBUF[29]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[2]_inst 
       (.I(D_MEM_ADDR_OBUF[2]),
        .O(D_MEM_ADDR[2]));
  LUT6 #(
    .INIT(64'hFF10FFFFFF100000)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[2]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[2]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[2]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[2]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[2]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[2]));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_17_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_18_n_0 ),
        .I3(ALU_DIN2[2]),
        .I4(\D_MEM_ADDR_OBUF[10]_inst_i_12_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[2]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_11 
       (.I0(ALU_DIN1[18]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[2]),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_2 
       (.I0(ID_EX_Q[81]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[2]),
        .I3(ALU_DIN2[2]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_3 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[2]),
        .I4(ALU_DIN1[2]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5404)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[2]_inst_i_7_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_12_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[2]_inst_i_8_n_0 ),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h020202A2)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_10_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[2]_inst_i_9_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_6 
       (.I0(\alu/data0 [2]),
        .I1(ID_EX_Q[125]),
        .I2(\alu/data1 [2]),
        .I3(ID_EX_Q[123]),
        .I4(ID_EX_Q[122]),
        .I5(\alu/data2 [2]),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_13_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[2]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[1]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEFFFEF)) 
    \D_MEM_ADDR_OBUF[2]_inst_i_9 
       (.I0(ALU_DIN2[2]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(EX_RF_RD1[1]),
        .I3(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I4(ID_EX_Q[127]),
        .I5(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[2]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[30]_inst 
       (.I(D_MEM_ADDR_OBUF[30]),
        .O(D_MEM_ADDR[30]));
  LUT6 #(
    .INIT(64'hFFFFBBABAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[30]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[30]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[30]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[30]));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_10 
       (.I0(ID_EX_Q[118]),
        .I1(ID_EX_Q[117]),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_16_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_11 
       (.I0(ALU_DIN2[2]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(ALU_DIN1[30]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_12 
       (.I0(ALU_DIN2[5]),
        .I1(\D_MEM_ADDR_OBUF[30]_inst_i_17_n_0 ),
        .I2(ALU_DIN2[15]),
        .I3(ALU_DIN2[16]),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_18_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_19_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_13 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_30_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_31_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[30]_inst_i_20_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_33_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h000000E2E2E200E2)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_14 
       (.I0(EX_RF_RD1[31]),
        .I1(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I2(ID_EX_Q[157]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0100FF010100FE00)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_15 
       (.I0(ALU_DIN2[2]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[30]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_16 
       (.I0(ALU_DIN2[1]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEA)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_17 
       (.I0(ALU_DIN2[30]),
        .I1(ID_EX_Q[110]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[31]),
        .I4(ALU_DIN2[22]),
        .I5(ALU_DIN2[6]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_18 
       (.I0(ALU_DIN2[11]),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN2[21]),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_35_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_19 
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN2[19]),
        .I3(ALU_DIN2[27]),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_27_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[31]_inst_i_26_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_2 
       (.I0(\alu/data0 [30]),
        .I1(ID_EX_Q[125]),
        .I2(\alu/data1 [30]),
        .I3(ID_EX_Q[123]),
        .I4(ID_EX_Q[122]),
        .I5(\alu/data2 [30]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_20 
       (.I0(ALU_DIN1[15]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[7]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[23]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_20_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_3 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(\D_MEM_ADDR_OBUF[30]_inst_i_8_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT5 #(
    .INIT(32'hFE0E0EFE)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_4 
       (.I0(ID_EX_Q[116]),
        .I1(ID_EX_Q[117]),
        .I2(ID_EX_Q[118]),
        .I3(ALU_DIN2[30]),
        .I4(ALU_DIN1[30]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3232320202020202)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[30]_inst_i_9_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[30]_inst_i_10_n_0 ),
        .I2(ID_EX_Q[117]),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_11_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h8A800000)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_6 
       (.I0(ID_EX_Q[121]),
        .I1(\D_MEM_ADDR_OBUF[30]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_10_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_7 
       (.I0(ID_EX_Q[123]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[125]),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_8 
       (.I0(ID_EX_Q[109]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[30]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFB80000)) 
    \D_MEM_ADDR_OBUF[30]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[30]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[30]_inst_i_15_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(ID_EX_Q[116]),
        .I5(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[30]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[31]_inst 
       (.I(D_MEM_ADDR_OBUF[31]),
        .O(D_MEM_ADDR[31]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAFE)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[31]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_4_n_0 ),
        .I3(ID_EX_Q[123]),
        .I4(ID_EX_Q[122]),
        .I5(ID_EX_Q[125]),
        .O(D_MEM_ADDR_OBUF[31]));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_22_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_23_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_24_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[31]_inst_i_25_n_0 ),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_11 
       (.I0(ID_EX_Q[121]),
        .I1(\D_MEM_ADDR_OBUF[31]_inst_i_26_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_27_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_28_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_29_n_0 ),
        .I5(ALU_DIN2[5]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h474747470033CCFF)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_30_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_31_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_32_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_33_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_13 
       (.I0(EX_RF_RD2[31]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[110]),
        .I3(EX_RF_RD1[31]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I5(ID_EX_Q[157]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_14 
       (.I0(EX_RF_RD2[30]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[109]),
        .I3(EX_RF_RD1[30]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I5(ID_EX_Q[156]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_15 
       (.I0(EX_RF_RD2[29]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[108]),
        .I3(EX_RF_RD1[29]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[155]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_16 
       (.I0(EX_RF_RD2[28]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[107]),
        .I3(EX_RF_RD1[28]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[154]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_17 
       (.I0(ID_EX_Q[157]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[31]),
        .I3(ID_EX_Q[110]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[31]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_18 
       (.I0(ID_EX_Q[156]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[30]),
        .I3(ID_EX_Q[109]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[30]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_19 
       (.I0(ID_EX_Q[155]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[29]),
        .I3(ID_EX_Q[108]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[29]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_2 
       (.I0(\alu/data0 [31]),
        .I1(ID_EX_Q[125]),
        .I2(\alu/data1 [31]),
        .I3(ID_EX_Q[123]),
        .I4(\alu/data2 [31]),
        .I5(ID_EX_Q[122]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_20 
       (.I0(ID_EX_Q[154]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[28]),
        .I3(ID_EX_Q[107]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[28]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_21 
       (.I0(ALU_DIN2[0]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN2[4]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_22 
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN1[16]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[8]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[24]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_23 
       (.I0(ALU_DIN1[4]),
        .I1(ALU_DIN1[20]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[12]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[28]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_24 
       (.I0(ALU_DIN1[2]),
        .I1(ALU_DIN1[18]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[10]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[26]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_25 
       (.I0(ALU_DIN1[6]),
        .I1(ALU_DIN1[22]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[14]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[30]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEA)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_26 
       (.I0(ALU_DIN2[29]),
        .I1(ID_EX_Q[88]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[9]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN2[10]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEA)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_27 
       (.I0(ALU_DIN2[23]),
        .I1(ID_EX_Q[96]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[17]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN2[12]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEA)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_28 
       (.I0(ALU_DIN2[27]),
        .I1(ID_EX_Q[98]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[19]),
        .I4(ALU_DIN2[14]),
        .I5(ALU_DIN2[8]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_29 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_34_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[31]_inst_i_35_n_0 ),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN2[13]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN2[11]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002EE2)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_8_n_0 ),
        .I1(ID_EX_Q[118]),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[31]),
        .I4(\D_MEM_ADDR_OBUF[29]_inst_i_7_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[31]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_30 
       (.I0(ALU_DIN1[1]),
        .I1(ALU_DIN1[17]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[9]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[25]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_31 
       (.I0(ALU_DIN1[5]),
        .I1(ALU_DIN1[21]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[13]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[29]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_32 
       (.I0(ALU_DIN1[7]),
        .I1(ALU_DIN1[23]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[15]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(\Q[63]_i_1__1_n_0 ),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_33 
       (.I0(ALU_DIN1[3]),
        .I1(ALU_DIN1[19]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[11]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[27]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_34 
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN2[15]),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN2[22]),
        .I4(ALU_DIN2[31]),
        .I5(ALU_DIN2[30]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEA)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_35 
       (.I0(ALU_DIN2[20]),
        .I1(ID_EX_Q[86]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(EX_RF_RD2[7]),
        .I4(ALU_DIN2[25]),
        .I5(ALU_DIN2[18]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_35_n_0 ));
  LUT4 #(
    .INIT(16'h880C)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_10_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_4_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[31]_inst_i_5 
       (.CI(\D_MEM_ADDR_OBUF[28]_inst_i_6_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[31]_inst_i_5_n_2 ,\D_MEM_ADDR_OBUF[31]_inst_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/data0 [31:29]),
        .S({\<const0> ,ID_EX_Q[157:155]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[31]_inst_i_6 
       (.CI(\D_MEM_ADDR_OBUF[27]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[31]_inst_i_6_n_1 ,\D_MEM_ADDR_OBUF[31]_inst_i_6_n_2 ,\D_MEM_ADDR_OBUF[31]_inst_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,ALU_DIN1[30:28]}),
        .O(\alu/data1 [31:28]),
        .S({\D_MEM_ADDR_OBUF[31]_inst_i_13_n_0 ,\D_MEM_ADDR_OBUF[31]_inst_i_14_n_0 ,\D_MEM_ADDR_OBUF[31]_inst_i_15_n_0 ,\D_MEM_ADDR_OBUF[31]_inst_i_16_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[31]_inst_i_7 
       (.CI(\D_MEM_ADDR_OBUF[27]_inst_i_7_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[31]_inst_i_7_n_1 ,\D_MEM_ADDR_OBUF[31]_inst_i_7_n_2 ,\D_MEM_ADDR_OBUF[31]_inst_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,ALU_DIN1[30:28]}),
        .O(\alu/data2 [31:28]),
        .S({\D_MEM_ADDR_OBUF[31]_inst_i_17_n_0 ,\D_MEM_ADDR_OBUF[31]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[31]_inst_i_19_n_0 ,\D_MEM_ADDR_OBUF[31]_inst_i_20_n_0 }));
  LUT6 #(
    .INIT(64'h000500050455FFFF)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[26]_inst_i_9_n_0 ),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_21_n_0 ),
        .I4(ID_EX_Q[116]),
        .I5(ID_EX_Q[117]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000000F010D0D0D0)) 
    \D_MEM_ADDR_OBUF[31]_inst_i_9 
       (.I0(ID_EX_Q[110]),
        .I1(ID_EX_Q[114]),
        .I2(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .I3(ALU_DIN2[31]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(ID_EX_Q[115]),
        .O(\D_MEM_ADDR_OBUF[31]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[3]_inst 
       (.I(D_MEM_ADDR_OBUF[3]),
        .O(D_MEM_ADDR[3]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[3]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_10 
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN2[2]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[2]),
        .I5(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[7]_inst_i_25_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_30_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[9]_inst_i_17_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_15_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_19_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[5]_inst_i_10_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_31_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_13 
       (.I0(ID_EX_Q[82]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[3]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_14 
       (.I0(ID_EX_Q[129]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[3]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_15 
       (.I0(ID_EX_Q[128]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[2]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_16 
       (.I0(ID_EX_Q[127]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[1]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_17 
       (.I0(ID_EX_Q[126]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[0]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hB847)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_18 
       (.I0(ID_EX_Q[129]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[3]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hB847)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_19 
       (.I0(ID_EX_Q[128]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[2]),
        .I3(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_2 
       (.I0(\alu/data2 [3]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [3]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [3]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hB847)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_20 
       (.I0(ID_EX_Q[127]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[1]),
        .I3(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hB847)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_21 
       (.I0(ID_EX_Q[126]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[0]),
        .I3(ALU_DIN2[0]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_22 
       (.I0(ID_EX_Q[129]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[3]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_23 
       (.I0(ID_EX_Q[128]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[2]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_24 
       (.I0(ID_EX_Q[127]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[1]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_25 
       (.I0(ID_EX_Q[126]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[0]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_26 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I1(EX_RF_RD1[3]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(ID_EX_Q[129]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_27 
       (.I0(ALU_DIN2[2]),
        .I1(EX_RF_RD1[2]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(ID_EX_Q[128]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_28 
       (.I0(ALU_DIN2[1]),
        .I1(EX_RF_RD1[1]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(ID_EX_Q[127]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_29 
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(ALU_DIN2[0]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[3]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_30 
       (.I0(ALU_DIN1[27]),
        .I1(ALU_DIN1[11]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[19]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[3]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_31 
       (.I0(\D_MEM_ADDR_OBUF[7]_inst_i_26_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_20_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_32_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_32 
       (.I0(ALU_DIN1[19]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[3]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[4]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_13_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN1[3]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[3]_inst_i_7 
       (.I0(ID_EX_Q[82]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[3]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[3]_inst_i_7_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[3]_inst_i_8 
       (.CI(\<const0> ),
        .CO({\D_MEM_ADDR_OBUF[3]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[3]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[3]_inst_i_8_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\D_MEM_ADDR_OBUF[3]_inst_i_14_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_15_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_16_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_17_n_0 }),
        .O(\alu/data2 [3:0]),
        .S({\D_MEM_ADDR_OBUF[3]_inst_i_18_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_19_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_20_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_21_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[3]_inst_i_9 
       (.CI(\<const0> ),
        .CO({\D_MEM_ADDR_OBUF[3]_inst_i_9_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_9_n_1 ,\D_MEM_ADDR_OBUF[3]_inst_i_9_n_2 ,\D_MEM_ADDR_OBUF[3]_inst_i_9_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\D_MEM_ADDR_OBUF[3]_inst_i_22_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_23_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_24_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_25_n_0 }),
        .O(\alu/data1 [3:0]),
        .S({\D_MEM_ADDR_OBUF[3]_inst_i_26_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_27_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_28_n_0 ,\D_MEM_ADDR_OBUF[3]_inst_i_29_n_0 }));
  OBUF \D_MEM_ADDR_OBUF[4]_inst 
       (.I(D_MEM_ADDR_OBUF[4]),
        .O(D_MEM_ADDR[4]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[4]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[4]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[4]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_17_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_15_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[7]_inst_i_24_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[7]_inst_i_25_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[8]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_16_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[9]_inst_i_15_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[6]_inst_i_11_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_17_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_18_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[10]_inst_i_10_n_0 ),
        .I4(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_13 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_19_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_20_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[8]_inst_i_15_n_0 ),
        .I4(ALU_DIN2[2]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_13_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_14 
       (.I0(ID_EX_Q[128]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_15 
       (.I0(ALU_DIN1[29]),
        .I1(ALU_DIN1[13]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[21]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[5]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_16 
       (.I0(ALU_DIN1[28]),
        .I1(ALU_DIN1[12]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[20]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[4]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_17 
       (.I0(ALU_DIN1[30]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[14]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_18 
       (.I0(ALU_DIN1[22]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[6]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_19 
       (.I0(ALU_DIN1[28]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[12]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_2 
       (.I0(\alu/data2 [4]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [4]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [4]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_20 
       (.I0(ALU_DIN1[20]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[4]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_9_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[5]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[4]_inst_i_10_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FF4747)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[4]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[4]_inst_i_13_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[5]_inst_i_7_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[4]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_7 
       (.I0(ID_EX_Q[83]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[4]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_7_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[4]_inst_i_8 
       (.CI(\<const0> ),
        .CO({\D_MEM_ADDR_OBUF[4]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[4]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[4]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[4]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,ID_EX_Q[128],\<const0> }),
        .O(\alu/data0 [4:1]),
        .S({ID_EX_Q[130:129],\D_MEM_ADDR_OBUF[4]_inst_i_14_n_0 ,ID_EX_Q[127]}));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \D_MEM_ADDR_OBUF[4]_inst_i_9 
       (.I0(ALU_DIN1[1]),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN2[2]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[3]),
        .I5(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[4]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[5]_inst 
       (.I(D_MEM_ADDR_OBUF[5]),
        .O(D_MEM_ADDR[5]));
  LUT6 #(
    .INIT(64'hFF10FFFFFF100000)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[5]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[5]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[5]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[5]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[5]_inst_i_6_n_0 ),
        .O(D_MEM_ADDR_OBUF[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_17_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[5]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_11 
       (.I0(ALU_DIN1[21]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[5]),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_2 
       (.I0(ID_EX_Q[84]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[5]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_3 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[5]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4540)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[6]_inst_i_10_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[5]_inst_i_7_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[5]_inst_i_8_n_0 ),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h08000888)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_5 
       (.I0(ID_EX_Q[121]),
        .I1(\D_MEM_ADDR_OBUF[30]_inst_i_12_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[5]_inst_i_9_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[6]_inst_i_8_n_0 ),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_6 
       (.I0(\alu/data0 [5]),
        .I1(ID_EX_Q[125]),
        .I2(\alu/data1 [5]),
        .I3(ID_EX_Q[123]),
        .I4(ID_EX_Q[122]),
        .I5(\alu/data2 [5]),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_7 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_19_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[5]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[7]_inst_i_12_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[6]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEF0000)) 
    \D_MEM_ADDR_OBUF[5]_inst_i_9 
       (.I0(ALU_DIN2[2]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(ALU_DIN1[2]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN2[1]),
        .I5(\D_MEM_ADDR_OBUF[7]_inst_i_23_n_0 ),
        .O(\D_MEM_ADDR_OBUF[5]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[6]_inst 
       (.I(D_MEM_ADDR_OBUF[6]),
        .O(D_MEM_ADDR[6]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[6]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[6]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[6]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[6]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[6]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[6]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[6]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[12]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[8]_inst_i_15_n_0 ),
        .I3(ALU_DIN2[1]),
        .I4(\D_MEM_ADDR_OBUF[4]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_11 
       (.I0(ALU_DIN1[30]),
        .I1(ALU_DIN1[14]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[22]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[6]),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_2 
       (.I0(\alu/data2 [6]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [6]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [6]),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[6]_inst_i_8_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[7]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[7]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[6]_inst_i_9_n_0 ),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF470047FF)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[7]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[6]_inst_i_10_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[6]),
        .I4(ALU_DIN1[6]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_7 
       (.I0(ID_EX_Q[85]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[6]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEF0000)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_8 
       (.I0(ALU_DIN2[2]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(ALU_DIN1[3]),
        .I3(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I4(ALU_DIN2[1]),
        .I5(\D_MEM_ADDR_OBUF[8]_inst_i_12_n_0 ),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[6]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_15_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[6]_inst_i_11_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[8]_inst_i_13_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[8]_inst_i_14_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[6]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[7]_inst 
       (.I(D_MEM_ADDR_OBUF[7]),
        .O(D_MEM_ADDR[7]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[7]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[7]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[7]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[7]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[7]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[7]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[7]_inst_i_23_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[7]_inst_i_24_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[7]_inst_i_25_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[9]_inst_i_16_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[9]_inst_i_17_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_18_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[7]_inst_i_26_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_13 
       (.I0(ID_EX_Q[130]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[4]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_14 
       (.I0(ID_EX_Q[133]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[7]),
        .I3(ID_EX_Q[86]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[7]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_15 
       (.I0(ID_EX_Q[132]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[6]),
        .I3(ID_EX_Q[85]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[6]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_16 
       (.I0(ID_EX_Q[131]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[5]),
        .I3(ID_EX_Q[84]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(EX_RF_RD2[5]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hB847)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_17 
       (.I0(ID_EX_Q[130]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[4]),
        .I3(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_18 
       (.I0(ID_EX_Q[130]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[4]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_19 
       (.I0(EX_RF_RD2[7]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[86]),
        .I3(EX_RF_RD1[7]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[133]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_2 
       (.I0(\alu/data2 [7]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [7]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [7]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_20 
       (.I0(EX_RF_RD2[6]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[85]),
        .I3(EX_RF_RD1[6]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[132]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_21 
       (.I0(EX_RF_RD2[5]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[84]),
        .I3(EX_RF_RD1[5]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I5(ID_EX_Q[131]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_22 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(EX_RF_RD1[4]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[130]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_23 
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[2]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN1[4]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_24 
       (.I0(ALU_DIN1[19]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[27]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[11]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_25 
       (.I0(\Q[63]_i_1__1_n_0 ),
        .I1(ALU_DIN1[15]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[23]),
        .I4(op_a2_carry_i_9_n_0),
        .I5(ALU_DIN1[7]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_26 
       (.I0(ALU_DIN2[5]),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(op_a2_carry_i_9_n_0),
        .I3(ALU_DIN1[15]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[7]_inst_i_27_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_27 
       (.I0(ALU_DIN1[23]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[7]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[7]_inst_i_10_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[8]_inst_i_9_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[8]_inst_i_10_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[7]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FF4747)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[7]_inst_i_12_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[8]_inst_i_11_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[7]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[7]_inst_i_7 
       (.I0(ID_EX_Q[86]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[7]),
        .I3(ALU_DIN2[7]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[7]_inst_i_7_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[7]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[3]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[7]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[7]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[7]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({ALU_DIN1[7:5],\D_MEM_ADDR_OBUF[7]_inst_i_13_n_0 }),
        .O(\alu/data2 [7:4]),
        .S({\D_MEM_ADDR_OBUF[7]_inst_i_14_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_15_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_16_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_17_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[7]_inst_i_9 
       (.CI(\D_MEM_ADDR_OBUF[3]_inst_i_9_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[7]_inst_i_9_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_9_n_1 ,\D_MEM_ADDR_OBUF[7]_inst_i_9_n_2 ,\D_MEM_ADDR_OBUF[7]_inst_i_9_n_3 }),
        .CYINIT(\<const0> ),
        .DI({ALU_DIN1[7:5],\D_MEM_ADDR_OBUF[7]_inst_i_18_n_0 }),
        .O(\alu/data1 [7:4]),
        .S({\D_MEM_ADDR_OBUF[7]_inst_i_19_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_20_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_21_n_0 ,\D_MEM_ADDR_OBUF[7]_inst_i_22_n_0 }));
  OBUF \D_MEM_ADDR_OBUF[8]_inst 
       (.I(D_MEM_ADDR_OBUF[8]),
        .O(D_MEM_ADDR[8]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[8]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[8]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[8]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[8]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[8]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[8]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_15_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[8]_inst_i_13_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[8]_inst_i_14_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[14]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[10]_inst_i_10_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[12]_inst_i_14_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[8]_inst_i_15_n_0 ),
        .I5(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_12 
       (.I0(ALU_DIN1[1]),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[5]),
        .I4(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_13 
       (.I0(ALU_DIN1[20]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[28]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[12]),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_14 
       (.I0(ALU_DIN1[16]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[24]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[8]),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4D48FFFF4D480000)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_15 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[16]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[8]_inst_i_16_n_0 ),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_16 
       (.I0(ALU_DIN1[24]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[8]),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_2 
       (.I0(\alu/data2 [8]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [8]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [8]),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[8]_inst_i_9_n_0 ),
        .I1(ALU_DIN2[0]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_8_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[9]_inst_i_10_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[8]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF470047FF)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_12_n_0 ),
        .I3(ALU_DIN2[0]),
        .I4(\D_MEM_ADDR_OBUF[8]_inst_i_11_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[8]),
        .I4(ALU_DIN1[8]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_7 
       (.I0(ID_EX_Q[87]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[8]),
        .I3(ALU_DIN2[8]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_7_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \D_MEM_ADDR_OBUF[8]_inst_i_8 
       (.CI(\D_MEM_ADDR_OBUF[4]_inst_i_8_n_0 ),
        .CO({\D_MEM_ADDR_OBUF[8]_inst_i_8_n_0 ,\D_MEM_ADDR_OBUF[8]_inst_i_8_n_1 ,\D_MEM_ADDR_OBUF[8]_inst_i_8_n_2 ,\D_MEM_ADDR_OBUF[8]_inst_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/data0 [8:5]),
        .S(ID_EX_Q[134:131]));
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[8]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[8]_inst_i_12_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[10]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[8]_inst_i_9_n_0 ));
  OBUF \D_MEM_ADDR_OBUF[9]_inst 
       (.I(D_MEM_ADDR_OBUF[9]),
        .O(D_MEM_ADDR[9]));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_1 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_2_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[9]_inst_i_3_n_0 ),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_4_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[9]_inst_i_5_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[9]_inst_i_6_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[9]_inst_i_7_n_0 ),
        .O(D_MEM_ADDR_OBUF[9]));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_10 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_16_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_17_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[11]_inst_i_22_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_11 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_15_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_18_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_12 
       (.I0(\D_MEM_ADDR_OBUF[13]_inst_i_16_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_19_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_13 
       (.I0(ALU_DIN1[2]),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I3(ALU_DIN1[6]),
        .I4(op_a2_carry_i_9_n_0),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_14 
       (.I0(ALU_DIN1[22]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[30]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[14]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_15 
       (.I0(ALU_DIN1[18]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[26]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[10]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_16 
       (.I0(ALU_DIN1[21]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[29]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[13]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_17 
       (.I0(ALU_DIN1[17]),
        .I1(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I2(ALU_DIN1[25]),
        .I3(op_a2_carry_i_9_n_0),
        .I4(ALU_DIN1[9]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h4D48FFFF4D480000)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_18 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[19]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[9]_inst_i_20_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4D48FFFF4D480000)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_19 
       (.I0(op_a2_carry_i_9_n_0),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[17]),
        .I4(\D_MEM_ADDR_OBUF[3]_inst_i_13_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[9]_inst_i_21_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_2 
       (.I0(\alu/data2 [9]),
        .I1(ID_EX_Q[122]),
        .I2(ID_EX_Q[123]),
        .I3(\alu/data1 [9]),
        .I4(ID_EX_Q[125]),
        .I5(\alu/data0 [9]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_20 
       (.I0(ALU_DIN1[27]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[11]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_21 
       (.I0(ALU_DIN1[25]),
        .I1(op_a2_carry_i_9_n_0),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[9]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h2A20FFFF)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_3 
       (.I0(\D_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[9]_inst_i_8_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[10]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEAEEAAA)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_4 
       (.I0(\D_MEM_ADDR_OBUF[28]_inst_i_8_n_0 ),
        .I1(\D_MEM_ADDR_OBUF[15]_inst_i_13_n_0 ),
        .I2(ALU_DIN2[0]),
        .I3(\D_MEM_ADDR_OBUF[9]_inst_i_9_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[9]_inst_i_10_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FF4747)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_5 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_11_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_12_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[10]_inst_i_7_n_0 ),
        .I4(ALU_DIN2[0]),
        .I5(\D_MEM_ADDR_OBUF[15]_inst_i_11_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFFFEFEFEFE)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_6 
       (.I0(ID_EX_Q[119]),
        .I1(ID_EX_Q[120]),
        .I2(ID_EX_Q[121]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN1[9]),
        .I5(ID_EX_Q[118]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000F1DDD00000000)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_7 
       (.I0(ID_EX_Q[88]),
        .I1(ID_EX_Q[114]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[9]),
        .I4(ID_EX_Q[115]),
        .I5(\D_MEM_ADDR_OBUF[29]_inst_i_13_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'h8B)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_8 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_13_n_0 ),
        .I1(ALU_DIN2[1]),
        .I2(\D_MEM_ADDR_OBUF[11]_inst_i_21_n_0 ),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \D_MEM_ADDR_OBUF[9]_inst_i_9 
       (.I0(\D_MEM_ADDR_OBUF[9]_inst_i_14_n_0 ),
        .I1(ALU_DIN2[2]),
        .I2(\D_MEM_ADDR_OBUF[9]_inst_i_15_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[12]_inst_i_13_n_0 ),
        .I4(ALU_DIN2[1]),
        .O(\D_MEM_ADDR_OBUF[9]_inst_i_9_n_0 ));
  OBUF \D_MEM_BE_OBUF[0]_inst 
       (.I(D_MEM_BE_OBUF[0]),
        .O(D_MEM_BE[0]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \D_MEM_BE_OBUF[0]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .O(D_MEM_BE_OBUF[0]));
  OBUF \D_MEM_BE_OBUF[1]_inst 
       (.I(D_MEM_BE_OBUF[1]),
        .O(D_MEM_BE[1]));
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT4 #(
    .INIT(16'h3332)) 
    \D_MEM_BE_OBUF[1]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(ID_EX_Q[161]),
        .I3(ID_EX_Q[160]),
        .O(D_MEM_BE_OBUF[1]));
  OBUF \D_MEM_BE_OBUF[2]_inst 
       (.I(D_MEM_BE_OBUF[2]),
        .O(D_MEM_BE[2]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT4 #(
    .INIT(16'h33F8)) 
    \D_MEM_BE_OBUF[2]_inst_i_1 
       (.I0(ID_EX_Q[161]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(ID_EX_Q[160]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .O(D_MEM_BE_OBUF[2]));
  OBUF \D_MEM_BE_OBUF[3]_inst 
       (.I(D_MEM_BE_OBUF[3]),
        .O(D_MEM_BE[3]));
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT4 #(
    .INIT(16'hFEF0)) 
    \D_MEM_BE_OBUF[3]_inst_i_1 
       (.I0(ID_EX_Q[161]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(ID_EX_Q[160]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .O(D_MEM_BE_OBUF[3]));
  OBUF D_MEM_CSN_OBUF_inst
       (.I(D_MEM_CSN_OBUF),
        .O(D_MEM_CSN));
  OBUF \D_MEM_DI_OBUF[0]_inst 
       (.I(D_MEM_DI_OBUF[0]),
        .O(D_MEM_DI[0]));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[0]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[0]),
        .O(D_MEM_DI_OBUF[0]));
  OBUF \D_MEM_DI_OBUF[10]_inst 
       (.I(D_MEM_DI_OBUF[10]),
        .O(D_MEM_DI[10]));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[10]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[2]),
        .I3(EX_RF_RD2[10]),
        .O(D_MEM_DI_OBUF[10]));
  OBUF \D_MEM_DI_OBUF[11]_inst 
       (.I(D_MEM_DI_OBUF[11]),
        .O(D_MEM_DI[11]));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[11]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[3]),
        .I3(EX_RF_RD2[11]),
        .O(D_MEM_DI_OBUF[11]));
  OBUF \D_MEM_DI_OBUF[12]_inst 
       (.I(D_MEM_DI_OBUF[12]),
        .O(D_MEM_DI[12]));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[12]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[4]),
        .I3(EX_RF_RD2[12]),
        .O(D_MEM_DI_OBUF[12]));
  OBUF \D_MEM_DI_OBUF[13]_inst 
       (.I(D_MEM_DI_OBUF[13]),
        .O(D_MEM_DI[13]));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[13]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[5]),
        .I3(EX_RF_RD2[13]),
        .O(D_MEM_DI_OBUF[13]));
  OBUF \D_MEM_DI_OBUF[14]_inst 
       (.I(D_MEM_DI_OBUF[14]),
        .O(D_MEM_DI[14]));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[14]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[6]),
        .I3(EX_RF_RD2[14]),
        .O(D_MEM_DI_OBUF[14]));
  OBUF \D_MEM_DI_OBUF[15]_inst 
       (.I(D_MEM_DI_OBUF[15]),
        .O(D_MEM_DI[15]));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[15]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[7]),
        .I3(EX_RF_RD2[15]),
        .O(D_MEM_DI_OBUF[15]));
  OBUF \D_MEM_DI_OBUF[16]_inst 
       (.I(D_MEM_DI_OBUF[16]),
        .O(D_MEM_DI[16]));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[16]_inst_i_1 
       (.I0(EX_RF_RD2[8]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[0]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[16]),
        .O(D_MEM_DI_OBUF[16]));
  OBUF \D_MEM_DI_OBUF[17]_inst 
       (.I(D_MEM_DI_OBUF[17]),
        .O(D_MEM_DI[17]));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[17]_inst_i_1 
       (.I0(EX_RF_RD2[9]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[1]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[17]),
        .O(D_MEM_DI_OBUF[17]));
  OBUF \D_MEM_DI_OBUF[18]_inst 
       (.I(D_MEM_DI_OBUF[18]),
        .O(D_MEM_DI[18]));
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[18]_inst_i_1 
       (.I0(EX_RF_RD2[10]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[2]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[18]),
        .O(D_MEM_DI_OBUF[18]));
  OBUF \D_MEM_DI_OBUF[19]_inst 
       (.I(D_MEM_DI_OBUF[19]),
        .O(D_MEM_DI[19]));
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[19]_inst_i_1 
       (.I0(EX_RF_RD2[11]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[3]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[19]),
        .O(D_MEM_DI_OBUF[19]));
  OBUF \D_MEM_DI_OBUF[1]_inst 
       (.I(D_MEM_DI_OBUF[1]),
        .O(D_MEM_DI[1]));
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[1]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[1]),
        .O(D_MEM_DI_OBUF[1]));
  OBUF \D_MEM_DI_OBUF[20]_inst 
       (.I(D_MEM_DI_OBUF[20]),
        .O(D_MEM_DI[20]));
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[20]_inst_i_1 
       (.I0(EX_RF_RD2[12]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[4]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[20]),
        .O(D_MEM_DI_OBUF[20]));
  OBUF \D_MEM_DI_OBUF[21]_inst 
       (.I(D_MEM_DI_OBUF[21]),
        .O(D_MEM_DI[21]));
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[21]_inst_i_1 
       (.I0(EX_RF_RD2[13]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[5]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[21]),
        .O(D_MEM_DI_OBUF[21]));
  OBUF \D_MEM_DI_OBUF[22]_inst 
       (.I(D_MEM_DI_OBUF[22]),
        .O(D_MEM_DI[22]));
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[22]_inst_i_1 
       (.I0(EX_RF_RD2[14]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[6]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[22]),
        .O(D_MEM_DI_OBUF[22]));
  OBUF \D_MEM_DI_OBUF[23]_inst 
       (.I(D_MEM_DI_OBUF[23]),
        .O(D_MEM_DI[23]));
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \D_MEM_DI_OBUF[23]_inst_i_1 
       (.I0(EX_RF_RD2[15]),
        .I1(D_MEM_ADDR_OBUF[0]),
        .I2(EX_RF_RD2[7]),
        .I3(D_MEM_ADDR_OBUF[1]),
        .I4(EX_RF_RD2[23]),
        .O(D_MEM_DI_OBUF[23]));
  OBUF \D_MEM_DI_OBUF[24]_inst 
       (.I(D_MEM_DI_OBUF[24]),
        .O(D_MEM_DI[24]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[24]_inst_i_1 
       (.I0(EX_RF_RD2[24]),
        .I1(EX_RF_RD2[8]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[0]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[16]),
        .O(D_MEM_DI_OBUF[24]));
  OBUF \D_MEM_DI_OBUF[25]_inst 
       (.I(D_MEM_DI_OBUF[25]),
        .O(D_MEM_DI[25]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[25]_inst_i_1 
       (.I0(EX_RF_RD2[25]),
        .I1(EX_RF_RD2[9]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[1]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[17]),
        .O(D_MEM_DI_OBUF[25]));
  OBUF \D_MEM_DI_OBUF[26]_inst 
       (.I(D_MEM_DI_OBUF[26]),
        .O(D_MEM_DI[26]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[26]_inst_i_1 
       (.I0(EX_RF_RD2[26]),
        .I1(EX_RF_RD2[10]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[2]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[18]),
        .O(D_MEM_DI_OBUF[26]));
  OBUF \D_MEM_DI_OBUF[27]_inst 
       (.I(D_MEM_DI_OBUF[27]),
        .O(D_MEM_DI[27]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[27]_inst_i_1 
       (.I0(EX_RF_RD2[27]),
        .I1(EX_RF_RD2[11]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[3]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[19]),
        .O(D_MEM_DI_OBUF[27]));
  OBUF \D_MEM_DI_OBUF[28]_inst 
       (.I(D_MEM_DI_OBUF[28]),
        .O(D_MEM_DI[28]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[28]_inst_i_1 
       (.I0(EX_RF_RD2[28]),
        .I1(EX_RF_RD2[12]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[4]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[20]),
        .O(D_MEM_DI_OBUF[28]));
  OBUF \D_MEM_DI_OBUF[29]_inst 
       (.I(D_MEM_DI_OBUF[29]),
        .O(D_MEM_DI[29]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[29]_inst_i_1 
       (.I0(EX_RF_RD2[29]),
        .I1(EX_RF_RD2[13]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[5]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[21]),
        .O(D_MEM_DI_OBUF[29]));
  OBUF \D_MEM_DI_OBUF[2]_inst 
       (.I(D_MEM_DI_OBUF[2]),
        .O(D_MEM_DI[2]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[2]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[2]),
        .O(D_MEM_DI_OBUF[2]));
  OBUF \D_MEM_DI_OBUF[30]_inst 
       (.I(D_MEM_DI_OBUF[30]),
        .O(D_MEM_DI[30]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[30]_inst_i_1 
       (.I0(EX_RF_RD2[30]),
        .I1(EX_RF_RD2[14]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[6]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[22]),
        .O(D_MEM_DI_OBUF[30]));
  OBUF \D_MEM_DI_OBUF[31]_inst 
       (.I(D_MEM_DI_OBUF[31]),
        .O(D_MEM_DI[31]));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \D_MEM_DI_OBUF[31]_inst_i_1 
       (.I0(EX_RF_RD2[31]),
        .I1(EX_RF_RD2[15]),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(EX_RF_RD2[7]),
        .I4(D_MEM_ADDR_OBUF[1]),
        .I5(EX_RF_RD2[23]),
        .O(D_MEM_DI_OBUF[31]));
  OBUF \D_MEM_DI_OBUF[3]_inst 
       (.I(D_MEM_DI_OBUF[3]),
        .O(D_MEM_DI[3]));
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[3]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[3]),
        .O(D_MEM_DI_OBUF[3]));
  OBUF \D_MEM_DI_OBUF[4]_inst 
       (.I(D_MEM_DI_OBUF[4]),
        .O(D_MEM_DI[4]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[4]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[4]),
        .O(D_MEM_DI_OBUF[4]));
  OBUF \D_MEM_DI_OBUF[5]_inst 
       (.I(D_MEM_DI_OBUF[5]),
        .O(D_MEM_DI[5]));
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[5]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[5]),
        .O(D_MEM_DI_OBUF[5]));
  OBUF \D_MEM_DI_OBUF[6]_inst 
       (.I(D_MEM_DI_OBUF[6]),
        .O(D_MEM_DI[6]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[6]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[6]),
        .O(D_MEM_DI_OBUF[6]));
  OBUF \D_MEM_DI_OBUF[7]_inst 
       (.I(D_MEM_DI_OBUF[7]),
        .O(D_MEM_DI[7]));
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \D_MEM_DI_OBUF[7]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[7]),
        .O(D_MEM_DI_OBUF[7]));
  OBUF \D_MEM_DI_OBUF[8]_inst 
       (.I(D_MEM_DI_OBUF[8]),
        .O(D_MEM_DI[8]));
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[8]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[0]),
        .I3(EX_RF_RD2[8]),
        .O(D_MEM_DI_OBUF[8]));
  OBUF \D_MEM_DI_OBUF[9]_inst 
       (.I(D_MEM_DI_OBUF[9]),
        .O(D_MEM_DI[9]));
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT4 #(
    .INIT(16'h3120)) 
    \D_MEM_DI_OBUF[9]_inst_i_1 
       (.I0(D_MEM_ADDR_OBUF[0]),
        .I1(D_MEM_ADDR_OBUF[1]),
        .I2(EX_RF_RD2[1]),
        .I3(EX_RF_RD2[9]),
        .O(D_MEM_DI_OBUF[9]));
  IBUF \D_MEM_DOUT_IBUF[0]_inst 
       (.I(D_MEM_DOUT[0]),
        .O(D_MEM_DOUT_IBUF[0]));
  IBUF \D_MEM_DOUT_IBUF[10]_inst 
       (.I(D_MEM_DOUT[10]),
        .O(D_MEM_DOUT_IBUF[10]));
  IBUF \D_MEM_DOUT_IBUF[11]_inst 
       (.I(D_MEM_DOUT[11]),
        .O(D_MEM_DOUT_IBUF[11]));
  IBUF \D_MEM_DOUT_IBUF[12]_inst 
       (.I(D_MEM_DOUT[12]),
        .O(D_MEM_DOUT_IBUF[12]));
  IBUF \D_MEM_DOUT_IBUF[13]_inst 
       (.I(D_MEM_DOUT[13]),
        .O(D_MEM_DOUT_IBUF[13]));
  IBUF \D_MEM_DOUT_IBUF[14]_inst 
       (.I(D_MEM_DOUT[14]),
        .O(D_MEM_DOUT_IBUF[14]));
  IBUF \D_MEM_DOUT_IBUF[15]_inst 
       (.I(D_MEM_DOUT[15]),
        .O(D_MEM_DOUT_IBUF[15]));
  IBUF \D_MEM_DOUT_IBUF[16]_inst 
       (.I(D_MEM_DOUT[16]),
        .O(D_MEM_DOUT_IBUF[16]));
  IBUF \D_MEM_DOUT_IBUF[17]_inst 
       (.I(D_MEM_DOUT[17]),
        .O(D_MEM_DOUT_IBUF[17]));
  IBUF \D_MEM_DOUT_IBUF[18]_inst 
       (.I(D_MEM_DOUT[18]),
        .O(D_MEM_DOUT_IBUF[18]));
  IBUF \D_MEM_DOUT_IBUF[19]_inst 
       (.I(D_MEM_DOUT[19]),
        .O(D_MEM_DOUT_IBUF[19]));
  IBUF \D_MEM_DOUT_IBUF[1]_inst 
       (.I(D_MEM_DOUT[1]),
        .O(D_MEM_DOUT_IBUF[1]));
  IBUF \D_MEM_DOUT_IBUF[20]_inst 
       (.I(D_MEM_DOUT[20]),
        .O(D_MEM_DOUT_IBUF[20]));
  IBUF \D_MEM_DOUT_IBUF[21]_inst 
       (.I(D_MEM_DOUT[21]),
        .O(D_MEM_DOUT_IBUF[21]));
  IBUF \D_MEM_DOUT_IBUF[22]_inst 
       (.I(D_MEM_DOUT[22]),
        .O(D_MEM_DOUT_IBUF[22]));
  IBUF \D_MEM_DOUT_IBUF[23]_inst 
       (.I(D_MEM_DOUT[23]),
        .O(D_MEM_DOUT_IBUF[23]));
  IBUF \D_MEM_DOUT_IBUF[24]_inst 
       (.I(D_MEM_DOUT[24]),
        .O(D_MEM_DOUT_IBUF[24]));
  IBUF \D_MEM_DOUT_IBUF[25]_inst 
       (.I(D_MEM_DOUT[25]),
        .O(D_MEM_DOUT_IBUF[25]));
  IBUF \D_MEM_DOUT_IBUF[26]_inst 
       (.I(D_MEM_DOUT[26]),
        .O(D_MEM_DOUT_IBUF[26]));
  IBUF \D_MEM_DOUT_IBUF[27]_inst 
       (.I(D_MEM_DOUT[27]),
        .O(D_MEM_DOUT_IBUF[27]));
  IBUF \D_MEM_DOUT_IBUF[28]_inst 
       (.I(D_MEM_DOUT[28]),
        .O(D_MEM_DOUT_IBUF[28]));
  IBUF \D_MEM_DOUT_IBUF[29]_inst 
       (.I(D_MEM_DOUT[29]),
        .O(D_MEM_DOUT_IBUF[29]));
  IBUF \D_MEM_DOUT_IBUF[2]_inst 
       (.I(D_MEM_DOUT[2]),
        .O(D_MEM_DOUT_IBUF[2]));
  IBUF \D_MEM_DOUT_IBUF[30]_inst 
       (.I(D_MEM_DOUT[30]),
        .O(D_MEM_DOUT_IBUF[30]));
  IBUF \D_MEM_DOUT_IBUF[31]_inst 
       (.I(D_MEM_DOUT[31]),
        .O(D_MEM_DOUT_IBUF[31]));
  IBUF \D_MEM_DOUT_IBUF[3]_inst 
       (.I(D_MEM_DOUT[3]),
        .O(D_MEM_DOUT_IBUF[3]));
  IBUF \D_MEM_DOUT_IBUF[4]_inst 
       (.I(D_MEM_DOUT[4]),
        .O(D_MEM_DOUT_IBUF[4]));
  IBUF \D_MEM_DOUT_IBUF[5]_inst 
       (.I(D_MEM_DOUT[5]),
        .O(D_MEM_DOUT_IBUF[5]));
  IBUF \D_MEM_DOUT_IBUF[6]_inst 
       (.I(D_MEM_DOUT[6]),
        .O(D_MEM_DOUT_IBUF[6]));
  IBUF \D_MEM_DOUT_IBUF[7]_inst 
       (.I(D_MEM_DOUT[7]),
        .O(D_MEM_DOUT_IBUF[7]));
  IBUF \D_MEM_DOUT_IBUF[8]_inst 
       (.I(D_MEM_DOUT[8]),
        .O(D_MEM_DOUT_IBUF[8]));
  IBUF \D_MEM_DOUT_IBUF[9]_inst 
       (.I(D_MEM_DOUT[9]),
        .O(D_MEM_DOUT_IBUF[9]));
  OBUF D_MEM_WEN_OBUF_inst
       (.I(D_MEM_WEN_OBUF),
        .O(D_MEM_WEN));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT2 #(
    .INIT(4'h8)) 
    D_MEM_WEN_OBUF_inst_i_1
       (.I0(ID_EX_Q[124]),
        .I1(RSTn_IBUF),
        .O(D_MEM_WEN_OBUF));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_ALU_SEL/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_ALU_SEL[26]),
        .Q(EX_CUSTOM_ALU_SEL[26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_ALU_SEL/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_ALU_SEL[27]),
        .Q(EX_CUSTOM_ALU_SEL[27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_ALU_SEL/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_ALU_SEL[28]),
        .Q(EX_CUSTOM_ALU_SEL[28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_ALU_SEL/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_ALU_SEL[29]),
        .Q(EX_CUSTOM_ALU_SEL[29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_ALU_SEL/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_ALU_SEL[30]),
        .Q(EX_CUSTOM_ALU_SEL[30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_ALU_SEL/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_ALU_SEL[31]),
        .Q(EX_CUSTOM_ALU_SEL[31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_EN/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_EN),
        .Q(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_RD/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(CUSTOM_RD),
        .Q(EX_CUSTOM_RD),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_RD_MEM/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(EX_CUSTOM_RD),
        .Q(MEM_CUSTOM_RD),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_CUSTOM_RD_WB/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(MEM_CUSTOM_RD),
        .Q(WB_CUSTOM_RD),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_Q[0]),
        .Q(EX_MEM_Q[0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[5]),
        .Q(EX_MEM_Q[10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[6]),
        .Q(EX_MEM_Q[11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[7]),
        .Q(EX_MEM_Q[12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[8]),
        .Q(EX_MEM_Q[13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[9]),
        .Q(EX_MEM_Q[14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[10]),
        .Q(EX_MEM_Q[15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[11]),
        .Q(EX_MEM_Q[16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[12]),
        .Q(EX_MEM_Q[17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[13]),
        .Q(EX_MEM_Q[18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[14]),
        .Q(EX_MEM_Q[19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_Q[1]),
        .Q(EX_MEM_Q[1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[15]),
        .Q(EX_MEM_Q[20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[16]),
        .Q(EX_MEM_Q[21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[17]),
        .Q(EX_MEM_Q[22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[18]),
        .Q(EX_MEM_Q[23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[19]),
        .Q(EX_MEM_Q[24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[20]),
        .Q(EX_MEM_Q[25]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[21]),
        .Q(EX_MEM_Q[26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[22]),
        .Q(EX_MEM_Q[27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[23]),
        .Q(EX_MEM_Q[28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[24]),
        .Q(EX_MEM_Q[29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_Q[2]),
        .Q(EX_MEM_Q[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[25]),
        .Q(EX_MEM_Q[30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[26]),
        .Q(EX_MEM_Q[31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[27]),
        .Q(EX_MEM_Q[32]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[28]),
        .Q(EX_MEM_Q[33]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[29]),
        .Q(EX_MEM_Q[34]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[30]),
        .Q(EX_MEM_Q[35]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[31]),
        .Q(EX_MEM_Q[36]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(D_MEM_CSN_OBUF),
        .Q(EX_MEM_Q[37]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_Q[113]),
        .Q(EX_MEM_Q[38]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_Q[124]),
        .Q(EX_MEM_Q[39]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_Q[3]),
        .Q(EX_MEM_Q[3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\FF_ID_EX/Q_reg_n_0_[164] ),
        .Q(MEM_LOAD_SEL[1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\FF_ID_EX/Q_reg_n_0_[165] ),
        .Q(MEM_LOAD_SEL[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\FF_ID_EX/Q_reg_n_0_[168] ),
        .Q(MEM_LOAD_SEL[5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\FF_ID_EX/Q_reg_n_0_[169] ),
        .Q(MEM_LOAD_SEL[6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_Q[4]),
        .Q(EX_MEM_Q[4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[0]),
        .Q(EX_MEM_Q[5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[1]),
        .Q(EX_MEM_Q[6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[2]),
        .Q(EX_MEM_Q[7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[3]),
        .Q(EX_MEM_Q[8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data0[4]),
        .Q(EX_MEM_Q[9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM_TEMP/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(D_MEM_ADDR_OBUF[0]),
        .Q(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_EX_MEM_TEMP/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(D_MEM_ADDR_OBUF[1]),
        .Q(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_DOUT_FILTERED[7]),
        .Q(ID_EX_Q[0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[100] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[21]),
        .Q(ID_EX_Q[100]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[101] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[22]),
        .Q(ID_EX_Q[101]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[102] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[23]),
        .Q(ID_EX_Q[102]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[103] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[24]),
        .Q(ID_EX_Q[103]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[104] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[25]),
        .Q(ID_EX_Q[104]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[105] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[26]),
        .Q(ID_EX_Q[105]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[106] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[27]),
        .Q(ID_EX_Q[106]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[107] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[28]),
        .Q(ID_EX_Q[107]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[108] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[29]),
        .Q(ID_EX_Q[108]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[109] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[30]),
        .Q(ID_EX_Q[109]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[110] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[31]),
        .Q(ID_EX_Q[110]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[112] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_D[112]),
        .Q(D_MEM_CSN_OBUF),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[113] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_WB_AFTER_LU),
        .Q(ID_EX_Q[113]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[114] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[20]),
        .Q(ID_EX_Q[114]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[115] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[21]),
        .Q(ID_EX_Q[115]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[116] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[22]),
        .Q(ID_EX_Q[116]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[117] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[23]),
        .Q(ID_EX_Q[117]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[118] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[24]),
        .Q(ID_EX_Q[118]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[119] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[25]),
        .Q(ID_EX_Q[119]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[120] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[26]),
        .Q(ID_EX_Q[120]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[121] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[27]),
        .Q(ID_EX_Q[121]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[122] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[28]),
        .Q(ID_EX_Q[122]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[123] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[29]),
        .Q(ID_EX_Q[123]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[124] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_D[124]),
        .Q(ID_EX_Q[124]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[125] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_JAL_AFTER_LU),
        .Q(ID_EX_Q[125]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[126] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[0]),
        .Q(ID_EX_Q[126]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[127] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[1]),
        .Q(ID_EX_Q[127]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[128] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[2]),
        .Q(ID_EX_Q[128]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[129] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[3]),
        .Q(ID_EX_Q[129]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[130] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[4]),
        .Q(ID_EX_Q[130]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[131] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[5]),
        .Q(ID_EX_Q[131]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[132] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[6]),
        .Q(ID_EX_Q[132]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[133] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[7]),
        .Q(ID_EX_Q[133]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[134] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[8]),
        .Q(ID_EX_Q[134]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[135] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[9]),
        .Q(ID_EX_Q[135]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[136] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[10]),
        .Q(ID_EX_Q[136]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[137] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[11]),
        .Q(ID_EX_Q[137]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[138] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[12]),
        .Q(ID_EX_Q[138]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[139] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[13]),
        .Q(ID_EX_Q[139]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[140] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[14]),
        .Q(ID_EX_Q[140]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[141] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[15]),
        .Q(ID_EX_Q[141]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[142] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[16]),
        .Q(ID_EX_Q[142]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[143] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[17]),
        .Q(ID_EX_Q[143]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[144] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[18]),
        .Q(ID_EX_Q[144]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[145] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[19]),
        .Q(ID_EX_Q[145]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[146] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[20]),
        .Q(ID_EX_Q[146]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[147] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[21]),
        .Q(ID_EX_Q[147]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[148] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[22]),
        .Q(ID_EX_Q[148]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[149] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[23]),
        .Q(ID_EX_Q[149]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[150] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[24]),
        .Q(ID_EX_Q[150]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[151] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[25]),
        .Q(ID_EX_Q[151]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[152] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[26]),
        .Q(ID_EX_Q[152]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[153] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[27]),
        .Q(ID_EX_Q[153]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[154] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[28]),
        .Q(ID_EX_Q[154]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[155] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[29]),
        .Q(ID_EX_Q[155]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[156] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[30]),
        .Q(ID_EX_Q[156]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[157] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_PC[31]),
        .Q(ID_EX_Q[157]),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[158]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[158] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE_EN),
        .Q(\FF_ID_EX/Q_reg_n_0_[158] ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[158]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[158]_rep 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[158]_rep_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[158]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[158]_rep__0 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[158]_rep__0_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[158]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[158]_rep__1 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[158]_rep__1_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[158]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[158]_rep__2 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[158]_rep__2_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[158]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[158]_rep__3 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[158]_rep__3_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[158]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[158]_rep__4 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[158]_rep__4_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[0]),
        .Q(EX_RF_RD2[0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[160] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[2]),
        .Q(ID_EX_Q[160]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[161] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[3]),
        .Q(ID_EX_Q[161]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[164] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[6]),
        .Q(\FF_ID_EX/Q_reg_n_0_[164] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[165] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[7]),
        .Q(\FF_ID_EX/Q_reg_n_0_[165] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[168] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[10]),
        .Q(\FF_ID_EX/Q_reg_n_0_[168] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[169] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[11]),
        .Q(\FF_ID_EX/Q_reg_n_0_[169] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[1]),
        .Q(EX_RF_RD2[1]),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[170]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[170] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[0]),
        .Q(\FF_ID_EX/Q_reg_n_0_[170] ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[170]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[170]_rep 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[170]_rep_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[170]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[170]_rep__0 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[170]_rep__0_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[170]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[170]_rep__1 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[170]_rep__1_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[170]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[170]_rep__2 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[170]_rep__2_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .R(RST0));
  (* ORIG_CELL_NAME = "Q_reg[170]" *) 
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[170]_rep__3 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[170]_rep__3_i_1_n_0 ),
        .Q(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[171] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_EX_D[171]),
        .Q(EX_BR_TAKEN),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[2]),
        .Q(EX_RF_RD2[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[3]),
        .Q(EX_RF_RD2[3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[4]),
        .Q(EX_RF_RD2[4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_DOUT_FILTERED[8]),
        .Q(ID_EX_Q[1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[5]),
        .Q(EX_RF_RD2[5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[6]),
        .Q(EX_RF_RD2[6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[7]),
        .Q(EX_RF_RD2[7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[8]),
        .Q(EX_RF_RD2[8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[9]),
        .Q(EX_RF_RD2[9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[10]),
        .Q(EX_RF_RD2[10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[11]),
        .Q(EX_RF_RD2[11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[12]),
        .Q(EX_RF_RD2[12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[13]),
        .Q(EX_RF_RD2[13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[14]),
        .Q(EX_RF_RD2[14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_DOUT_FILTERED[9]),
        .Q(ID_EX_Q[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[15]),
        .Q(EX_RF_RD2[15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[16]),
        .Q(EX_RF_RD2[16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[17]),
        .Q(EX_RF_RD2[17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[18]),
        .Q(EX_RF_RD2[18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[19]),
        .Q(EX_RF_RD2[19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[20]),
        .Q(EX_RF_RD2[20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[21]),
        .Q(EX_RF_RD2[21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[22]),
        .Q(EX_RF_RD2[22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[23]),
        .Q(EX_RF_RD2[23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[24]),
        .Q(EX_RF_RD2[24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_DOUT_FILTERED[10]),
        .Q(ID_EX_Q[3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[25]),
        .Q(EX_RF_RD2[25]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[26]),
        .Q(EX_RF_RD2[26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[27]),
        .Q(EX_RF_RD2[27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[28]),
        .Q(EX_RF_RD2[28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[29]),
        .Q(EX_RF_RD2[29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[30]),
        .Q(EX_RF_RD2[30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_RD2_FORWARDED[31]),
        .Q(EX_RF_RD2[31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[47]_i_1_n_0 ),
        .Q(EX_RF_RD1[0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[48]_i_1_n_0 ),
        .Q(EX_RF_RD1[1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[49] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[49]_i_1_n_0 ),
        .Q(EX_RF_RD1[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_DOUT_FILTERED[11]),
        .Q(ID_EX_Q[4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[50] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[50]_i_1_n_0 ),
        .Q(EX_RF_RD1[3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[51] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[51]_i_1_n_0 ),
        .Q(EX_RF_RD1[4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[52] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[52]_i_1_n_0 ),
        .Q(EX_RF_RD1[5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[53] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[53]_i_1_n_0 ),
        .Q(EX_RF_RD1[6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[54] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[54]_i_1_n_0 ),
        .Q(EX_RF_RD1[7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[55]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[56]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[57]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[58]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[59]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[60]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[61]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[62]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[63]_i_1_n_0 ),
        .Q(EX_RF_RD1[16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[64] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[64]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[65] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[65]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[66] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[66]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[67] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[67]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[68] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[68]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[69] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[69]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[70] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[70]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[71] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[71]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[72] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[72]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[25]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[73] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[73]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[74] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[74]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[75] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[75]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[76] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[76]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[77] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[77]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[78] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[78]_i_1__0_n_0 ),
        .Q(EX_RF_RD1[31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[79] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[0]),
        .Q(ID_EX_Q[79]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[80] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[1]),
        .Q(ID_EX_Q[80]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[81] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[2]),
        .Q(ID_EX_Q[81]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[82] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[3]),
        .Q(ID_EX_Q[82]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[83] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[4]),
        .Q(ID_EX_Q[83]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[84] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[5]),
        .Q(ID_EX_Q[84]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[85] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[6]),
        .Q(ID_EX_Q[85]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[86] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[7]),
        .Q(ID_EX_Q[86]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[87] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[8]),
        .Q(ID_EX_Q[87]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[88] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[9]),
        .Q(ID_EX_Q[88]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[89] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[10]),
        .Q(ID_EX_Q[89]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[90] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[11]),
        .Q(ID_EX_Q[90]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[91] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[12]),
        .Q(ID_EX_Q[91]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[92] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[13]),
        .Q(ID_EX_Q[92]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[93] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[14]),
        .Q(ID_EX_Q[93]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[94] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[15]),
        .Q(ID_EX_Q[94]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[95] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[16]),
        .Q(ID_EX_Q[95]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[96] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[17]),
        .Q(ID_EX_Q[96]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[97] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[18]),
        .Q(ID_EX_Q[97]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[98] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[19]),
        .Q(ID_EX_Q[98]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_ID_EX/Q_reg[99] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ID_IMMEDIATE[20]),
        .Q(ID_EX_Q[99]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[0]),
        .Q(ID_PC[0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[10]),
        .Q(ID_PC[10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[11]),
        .Q(ID_PC[11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[12]),
        .Q(ID_PC[12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[13]),
        .Q(ID_PC[13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[14]),
        .Q(ID_PC[14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[15]),
        .Q(ID_PC[15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[16]),
        .Q(ID_PC[16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[17]),
        .Q(ID_PC[17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[18]),
        .Q(ID_PC[18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[19]),
        .Q(ID_PC[19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[1]),
        .Q(ID_PC[1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[20]),
        .Q(ID_PC[20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[21]),
        .Q(ID_PC[21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[22]),
        .Q(ID_PC[22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[23]),
        .Q(ID_PC[23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[24]),
        .Q(ID_PC[24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[25]),
        .Q(ID_PC[25]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[26]),
        .Q(ID_PC[26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[27]),
        .Q(ID_PC[27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[28]),
        .Q(ID_PC[28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[29]),
        .Q(ID_PC[29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[2]),
        .Q(ID_PC[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[30]),
        .Q(ID_PC[30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[31]),
        .Q(ID_PC[31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[3]),
        .Q(ID_PC[3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[4]),
        .Q(ID_PC[4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[5]),
        .Q(ID_PC[5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[6]),
        .Q(ID_PC[6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[7]),
        .Q(ID_PC[7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[8]),
        .Q(ID_PC[8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PC/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(I_MEM_ADDR_OBUF[9]),
        .Q(ID_PC[9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[0]_i_1__4_n_0 ),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[10]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[11]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[12]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[13]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[14]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[15]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[16]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[17]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[18]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[19]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[1]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[20]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[21]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[22]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[23]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[24]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[25]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[26]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[27]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[28]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[29]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[2]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(D0),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[31]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[3]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[4]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[5]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[6]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[7]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[8]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_IF_ID_PCADD/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(IF_PC_ADD4[9]),
        .Q(\FF_IF_ID_PCADD/Q_reg_n_0_[9] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_JALR_EN/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(DECODED_INSTRUCTION[12]),
        .Q(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(EX_MEM_Q[0]),
        .Q(CRF_WA_OBUF[0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[5]),
        .Q(CRF_WD_OBUF[5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[6]),
        .Q(CRF_WD_OBUF[6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[7]),
        .Q(CRF_WD_OBUF[7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[8]),
        .Q(CRF_WD_OBUF[8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[9]),
        .Q(CRF_WD_OBUF[9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[10]),
        .Q(CRF_WD_OBUF[10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[11]),
        .Q(CRF_WD_OBUF[11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[12]),
        .Q(CRF_WD_OBUF[12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[13]),
        .Q(CRF_WD_OBUF[13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[14]),
        .Q(CRF_WD_OBUF[14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(EX_MEM_Q[1]),
        .Q(CRF_WA_OBUF[1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[15]),
        .Q(CRF_WD_OBUF[15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[16]),
        .Q(CRF_WD_OBUF[16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[17]),
        .Q(CRF_WD_OBUF[17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[18]),
        .Q(CRF_WD_OBUF[18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[19]),
        .Q(CRF_WD_OBUF[19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[20]),
        .Q(CRF_WD_OBUF[20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[21]),
        .Q(CRF_WD_OBUF[21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[22]),
        .Q(CRF_WD_OBUF[22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[23]),
        .Q(CRF_WD_OBUF[23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[24]),
        .Q(CRF_WD_OBUF[24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(EX_MEM_Q[2]),
        .Q(CRF_WA_OBUF[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[25]),
        .Q(CRF_WD_OBUF[25]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[26]),
        .Q(CRF_WD_OBUF[26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[27]),
        .Q(CRF_WD_OBUF[27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[28]),
        .Q(CRF_WD_OBUF[28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[29]),
        .Q(CRF_WD_OBUF[29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[30]),
        .Q(CRF_WD_OBUF[30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[31]),
        .Q(CRF_WD_OBUF[31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(EX_MEM_Q[38]),
        .Q(MEM_WB_Q),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(EX_MEM_Q[3]),
        .Q(CRF_WA_OBUF[3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(EX_MEM_Q[4]),
        .Q(CRF_WA_OBUF[4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[0]),
        .Q(CRF_WD_OBUF[0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[1]),
        .Q(CRF_WD_OBUF[1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[2]),
        .Q(CRF_WD_OBUF[2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[3]),
        .Q(CRF_WD_OBUF[3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_MEM_WB/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(data1[4]),
        .Q(CRF_WD_OBUF[4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[0]),
        .Q(STALL_COUNTER_Q[0]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[1]),
        .Q(STALL_COUNTER_Q[1]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[2]),
        .Q(STALL_COUNTER_Q[2]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[3]),
        .Q(STALL_COUNTER_Q[3]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[4]),
        .Q(STALL_COUNTER_Q[4]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[5]),
        .Q(STALL_COUNTER_Q[5]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[6]),
        .Q(STALL_COUNTER_Q[6]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[7]),
        .Q(STALL_COUNTER_Q[7]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[8]),
        .Q(STALL_COUNTER_Q[8]),
        .R(RST02_out));
  FDRE #(
    .INIT(1'b0)) 
    \FF_STALL_COUNTER/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(STALL_COUNTER_D[9]),
        .Q(STALL_COUNTER_Q[9]),
        .R(RST02_out));
  GND GND
       (.G(\<const0> ));
  GND GND_1
       (.G(GND_2));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__0_i_1
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__0_i_5_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__0_i_6_n_0),
        .O(\custom_alu/fp2int/p_0_in [8]));
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    INT0_carry__0_i_10
       (.I0(ALU_DIN1[18]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[10]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(INT0_carry__0_i_18_n_0),
        .I5(INT0_carry__0_i_21_n_0),
        .O(INT0_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    INT0_carry__0_i_11
       (.I0(ALU_DIN1[16]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[8]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(INT0_carry__0_i_18_n_0),
        .I5(INT0_carry__0_i_22_n_0),
        .O(INT0_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    INT0_carry__0_i_12
       (.I0(ALU_DIN1[19]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[11]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(INT0_carry__0_i_18_n_0),
        .I5(INT0_carry__0_i_23_n_0),
        .O(INT0_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    INT0_carry__0_i_13
       (.I0(ALU_DIN1[17]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[9]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(INT0_carry__0_i_18_n_0),
        .I5(INT0_carry__0_i_15_n_0),
        .O(INT0_carry__0_i_13_n_0));
  LUT6 #(
    .INIT(64'h44477747FFFFFFFF)) 
    INT0_carry__0_i_14
       (.I0(ALU_DIN1[17]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(EX_RF_RD1[9]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[135]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry__0_i_14_n_0));
  LUT6 #(
    .INIT(64'h44477747FFFFFFFF)) 
    INT0_carry__0_i_15
       (.I0(ALU_DIN1[21]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(EX_RF_RD1[13]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[139]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry__0_i_15_n_0));
  LUT5 #(
    .INIT(32'hCCA533A5)) 
    INT0_carry__0_i_16
       (.I0(EX_RF_RD1[23]),
        .I1(ID_EX_Q[149]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I4(ID_EX_Q[150]),
        .O(INT0_carry__0_i_16_n_0));
  LUT6 #(
    .INIT(64'h00FFFFFF47004700)) 
    INT0_carry__0_i_17
       (.I0(ID_EX_Q[133]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[7]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[15]),
        .I5(INT0_carry__2_i_13_n_0),
        .O(INT0_carry__0_i_17_n_0));
  LUT6 #(
    .INIT(64'h3C553CAACCAACCAA)) 
    INT0_carry__0_i_18
       (.I0(EX_RF_RD1[25]),
        .I1(ID_EX_Q[151]),
        .I2(ID_EX_Q[150]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[24]),
        .I5(ALU_DIN1[23]),
        .O(INT0_carry__0_i_18_n_0));
  LUT6 #(
    .INIT(64'h1D001DFFFFFFFFFF)) 
    INT0_carry__0_i_19
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(ALU_DIN1[11]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry__0_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__0_i_2
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__0_i_7_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__0_i_5_n_0),
        .O(\custom_alu/fp2int/p_0_in [7]));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__0_i_20
       (.I0(INT0_carry__0_i_11_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry_i_21_n_0),
        .O(INT0_carry__0_i_20_n_0));
  LUT6 #(
    .INIT(64'h44477747FFFFFFFF)) 
    INT0_carry__0_i_21
       (.I0(ALU_DIN1[22]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(EX_RF_RD1[14]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I4(ID_EX_Q[140]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry__0_i_21_n_0));
  LUT6 #(
    .INIT(64'h1D001DFFFFFFFFFF)) 
    INT0_carry__0_i_22
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(ALU_DIN1[12]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry__0_i_22_n_0));
  LUT6 #(
    .INIT(64'hDCCCCCCCC7777777)) 
    INT0_carry__0_i_23
       (.I0(ALU_DIN1[15]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN1[24]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN1[26]),
        .O(INT0_carry__0_i_23_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry__0_i_3
       (.I0(INT0_carry__0_i_8_n_0),
        .O(\custom_alu/fp2int/p_0_in [6]));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry__0_i_4
       (.I0(INT0_carry__0_i_9_n_0),
        .O(\custom_alu/fp2int/p_0_in [5]));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__0_i_5
       (.I0(INT0_carry__0_i_10_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__0_i_11_n_0),
        .O(INT0_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__0_i_6
       (.I0(INT0_carry__0_i_12_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__0_i_13_n_0),
        .O(INT0_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    INT0_carry__0_i_7
       (.I0(INT0_carry__0_i_14_n_0),
        .I1(INT0_carry__0_i_15_n_0),
        .I2(INT0_carry__0_i_16_n_0),
        .I3(INT0_carry__0_i_17_n_0),
        .I4(INT0_carry__0_i_18_n_0),
        .I5(INT0_carry__0_i_19_n_0),
        .O(INT0_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000101555551015)) 
    INT0_carry__0_i_8
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry_i_21_n_0),
        .I2(ALU_DIN1[24]),
        .I3(INT0_carry__0_i_11_n_0),
        .I4(ALU_DIN1[23]),
        .I5(INT0_carry__0_i_7_n_0),
        .O(INT0_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry__0_i_9
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry_i_10_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__0_i_20_n_0),
        .O(INT0_carry__0_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry__1_i_1
       (.I0(INT0_carry__1_i_5_n_0),
        .O(\custom_alu/fp2int/p_0_in [12]));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__1_i_10
       (.I0(INT0_carry__2_i_15_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__1_i_11_n_0),
        .O(INT0_carry__1_i_10_n_0));
  LUT6 #(
    .INIT(64'h5FFF30FF5FFF3FFF)) 
    INT0_carry__1_i_11
       (.I0(ALU_DIN1[21]),
        .I1(ALU_DIN1[13]),
        .I2(INT0_carry__0_i_18_n_0),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(INT0_carry__2_i_13_n_0),
        .I5(ALU_DIN1[17]),
        .O(INT0_carry__1_i_11_n_0));
  LUT6 #(
    .INIT(64'h5FFF30FF5FFF3FFF)) 
    INT0_carry__1_i_12
       (.I0(ALU_DIN1[22]),
        .I1(ALU_DIN1[14]),
        .I2(INT0_carry__0_i_18_n_0),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(INT0_carry__2_i_13_n_0),
        .I5(ALU_DIN1[18]),
        .O(INT0_carry__1_i_12_n_0));
  LUT6 #(
    .INIT(64'h5FFF30FF5FFF3FFF)) 
    INT0_carry__1_i_13
       (.I0(ALU_DIN1[20]),
        .I1(ALU_DIN1[12]),
        .I2(INT0_carry__0_i_18_n_0),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(INT0_carry__2_i_13_n_0),
        .I5(ALU_DIN1[16]),
        .O(INT0_carry__1_i_13_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__1_i_14
       (.I0(INT0_carry__1_i_13_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__0_i_10_n_0),
        .O(INT0_carry__1_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__1_i_2
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__1_i_6_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__1_i_7_n_0),
        .O(INT0_carry__1_i_2_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry__1_i_3
       (.I0(INT0_carry__1_i_8_n_0),
        .O(\custom_alu/fp2int/p_0_in [10]));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry__1_i_4
       (.I0(INT0_carry__1_i_9_n_0),
        .O(\custom_alu/fp2int/p_0_in [9]));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry__1_i_5
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__1_i_7_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__1_i_10_n_0),
        .O(INT0_carry__1_i_5_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__1_i_6
       (.I0(INT0_carry__1_i_11_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__0_i_12_n_0),
        .O(INT0_carry__1_i_6_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__1_i_7
       (.I0(INT0_carry__1_i_12_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__1_i_13_n_0),
        .O(INT0_carry__1_i_7_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry__1_i_8
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__1_i_14_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__1_i_6_n_0),
        .O(INT0_carry__1_i_8_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry__1_i_9
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__0_i_6_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__1_i_14_n_0),
        .O(INT0_carry__1_i_9_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__2_i_1
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__2_i_5_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__2_i_6_n_0),
        .O(INT0_carry__2_i_1_n_0));
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    INT0_carry__2_i_10
       (.I0(ALU_DIN1[18]),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(INT0_carry__2_i_13_n_0),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[22]),
        .O(INT0_carry__2_i_10_n_0));
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    INT0_carry__2_i_11
       (.I0(ALU_DIN1[16]),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(INT0_carry__2_i_13_n_0),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[20]),
        .O(INT0_carry__2_i_11_n_0));
  LUT5 #(
    .INIT(32'h55556AAA)) 
    INT0_carry__2_i_12
       (.I0(ALU_DIN1[27]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN1[24]),
        .I3(ALU_DIN1[23]),
        .I4(ALU_DIN1[26]),
        .O(INT0_carry__2_i_12_n_0));
  LUT6 #(
    .INIT(64'h1DE2E2E2E2E2E2E2)) 
    INT0_carry__2_i_13
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(ALU_DIN1[23]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN1[25]),
        .O(INT0_carry__2_i_13_n_0));
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    INT0_carry__2_i_14
       (.I0(ALU_DIN1[17]),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(INT0_carry__2_i_13_n_0),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[21]),
        .O(INT0_carry__2_i_14_n_0));
  LUT6 #(
    .INIT(64'h2F30AFFF2F3FAFFF)) 
    INT0_carry__2_i_15
       (.I0(ALU_DIN1[27]),
        .I1(ALU_DIN1[15]),
        .I2(INT0_carry__0_i_18_n_0),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(INT0_carry__2_i_12_n_0),
        .I5(ALU_DIN1[19]),
        .O(INT0_carry__2_i_15_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__2_i_16
       (.I0(INT0_carry__2_i_11_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__1_i_12_n_0),
        .O(INT0_carry__2_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__2_i_2
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__2_i_7_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__2_i_5_n_0),
        .O(INT0_carry__2_i_2_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry__2_i_3
       (.I0(INT0_carry__2_i_8_n_0),
        .O(\custom_alu/fp2int/p_0_in [14]));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry__2_i_4
       (.I0(INT0_carry__2_i_9_n_0),
        .O(\custom_alu/fp2int/p_0_in [13]));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__2_i_5
       (.I0(INT0_carry__2_i_10_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__2_i_11_n_0),
        .O(INT0_carry__2_i_5_n_0));
  LUT6 #(
    .INIT(64'hDFDDFFFFDFDD0000)) 
    INT0_carry__2_i_6
       (.I0(INT0_carry__2_i_12_n_0),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[19]),
        .I3(INT0_carry__0_i_18_n_0),
        .I4(INT0_carry__0_i_16_n_0),
        .I5(INT0_carry__2_i_14_n_0),
        .O(INT0_carry__2_i_6_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry__2_i_7
       (.I0(INT0_carry__2_i_14_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry__2_i_15_n_0),
        .O(INT0_carry__2_i_7_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry__2_i_8
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__2_i_16_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__2_i_7_n_0),
        .O(INT0_carry__2_i_8_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry__2_i_9
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__1_i_10_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__2_i_16_n_0),
        .O(INT0_carry__2_i_9_n_0));
  LUT6 #(
    .INIT(64'hFEFEAEAEFEFEAEFE)) 
    INT0_carry__3_i_1
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__3_i_5_n_0),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN1[24]),
        .I4(INT0_carry__3_i_6_n_0),
        .I5(ALU_DIN1[21]),
        .O(INT0_carry__3_i_1_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__3_i_2
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__3_i_7_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__3_i_5_n_0),
        .O(INT0_carry__3_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__3_i_3
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__3_i_8_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__3_i_7_n_0),
        .O(INT0_carry__3_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry__3_i_4
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__2_i_6_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__3_i_8_n_0),
        .O(INT0_carry__3_i_4_n_0));
  LUT6 #(
    .INIT(64'hFF4FFFFFFF7FFFFF)) 
    INT0_carry__3_i_5
       (.I0(ALU_DIN1[22]),
        .I1(INT0_carry__0_i_16_n_0),
        .I2(INT0_carry__0_i_18_n_0),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(INT0_carry__2_i_12_n_0),
        .I5(ALU_DIN1[20]),
        .O(INT0_carry__3_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT5 #(
    .INIT(32'hFDDDDFFF)) 
    INT0_carry__3_i_6
       (.I0(ALU_DIN1[27]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN1[24]),
        .I4(ALU_DIN1[25]),
        .O(INT0_carry__3_i_6_n_0));
  LUT6 #(
    .INIT(64'hFF4FFF7FFFCFFFCF)) 
    INT0_carry__3_i_7
       (.I0(ALU_DIN1[21]),
        .I1(INT0_carry__0_i_16_n_0),
        .I2(INT0_carry__2_i_12_n_0),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(ALU_DIN1[19]),
        .I5(INT0_carry__0_i_18_n_0),
        .O(INT0_carry__3_i_7_n_0));
  LUT6 #(
    .INIT(64'hDFFFFFFFDFFF0000)) 
    INT0_carry__3_i_8
       (.I0(INT0_carry__0_i_18_n_0),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(INT0_carry__2_i_12_n_0),
        .I3(ALU_DIN1[20]),
        .I4(INT0_carry__0_i_16_n_0),
        .I5(INT0_carry__2_i_10_n_0),
        .O(INT0_carry__3_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF77CF47)) 
    INT0_carry__4_i_1
       (.I0(ID_EX_Q[150]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[24]),
        .I3(ID_EX_Q[149]),
        .I4(EX_RF_RD1[23]),
        .I5(INT0_carry__4_i_4_n_0),
        .O(\custom_alu/fp2int/p_0_in [23]));
  LUT6 #(
    .INIT(64'hFFFFAAAAABFBFFFF)) 
    INT0_carry__4_i_2
       (.I0(INT0_carry__4_i_4_n_0),
        .I1(EX_RF_RD1[22]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(ID_EX_Q[148]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN1[23]),
        .O(INT0_carry__4_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFCFFF44)) 
    INT0_carry__4_i_3
       (.I0(ALU_DIN1[22]),
        .I1(ALU_DIN1[23]),
        .I2(ALU_DIN1[21]),
        .I3(INT0_carry__3_i_6_n_0),
        .I4(ALU_DIN1[24]),
        .I5(INT0_carry_i_6_n_0),
        .O(\custom_alu/fp2int/p_0_in [21]));
  LUT6 #(
    .INIT(64'hFFFFEBBBFFFFFFFF)) 
    INT0_carry__4_i_4
       (.I0(INT0_carry__4_i_5_n_0),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN1[24]),
        .I3(ALU_DIN1[23]),
        .I4(ALU_DIN1[26]),
        .I5(ALU_DIN1[27]),
        .O(INT0_carry__4_i_4_n_0));
  LUT6 #(
    .INIT(64'hBFFFFFFDFDFDFDFD)) 
    INT0_carry__4_i_5
       (.I0(ALU_DIN1[30]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN1[29]),
        .I3(INT0_carry__4_i_6_n_0),
        .I4(ALU_DIN1[26]),
        .I5(ALU_DIN1[27]),
        .O(INT0_carry__4_i_5_n_0));
  LUT6 #(
    .INIT(64'hC0AAC00000000000)) 
    INT0_carry__4_i_6
       (.I0(EX_RF_RD1[25]),
        .I1(ID_EX_Q[151]),
        .I2(ID_EX_Q[150]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[24]),
        .I5(ALU_DIN1[23]),
        .O(INT0_carry__4_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry_i_1
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry_i_7_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry_i_8_n_0),
        .O(\custom_alu/fp2int/p_0_in [0]));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry_i_10
       (.I0(INT0_carry_i_23_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry_i_24_n_0),
        .O(INT0_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry_i_11
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry_i_25_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry_i_9_n_0),
        .O(INT0_carry_i_11_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry_i_12
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry_i_26_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry_i_25_n_0),
        .O(INT0_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h0001110155511151)) 
    INT0_carry_i_13
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry_i_8_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry_i_26_n_0),
        .O(INT0_carry_i_13_n_0));
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT5 #(
    .INIT(32'hAAAA8000)) 
    INT0_carry_i_14
       (.I0(ALU_DIN1[27]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN1[24]),
        .I3(ALU_DIN1[23]),
        .I4(ALU_DIN1[26]),
        .O(INT0_carry_i_14_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    INT0_carry_i_15
       (.I0(INT0_carry_i_27_n_0),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(INT0_carry_i_28_n_0),
        .O(INT0_carry_i_15_n_0));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    INT0_carry_i_16
       (.I0(ALU_DIN1[8]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[0]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[16]),
        .O(INT0_carry_i_16_n_0));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    INT0_carry_i_17
       (.I0(ALU_DIN1[12]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[4]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[20]),
        .O(INT0_carry_i_17_n_0));
  LUT6 #(
    .INIT(64'h88BBBBBB8B888B88)) 
    INT0_carry_i_18
       (.I0(INT0_carry_i_29_n_0),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(ALU_DIN1[7]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[15]),
        .I5(INT0_carry__2_i_13_n_0),
        .O(INT0_carry_i_18_n_0));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    INT0_carry_i_19
       (.I0(ALU_DIN1[9]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[1]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[17]),
        .O(INT0_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    INT0_carry_i_2
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry_i_9_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry_i_10_n_0),
        .O(\custom_alu/fp2int/p_0_in [4]));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    INT0_carry_i_20
       (.I0(ALU_DIN1[13]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[5]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[21]),
        .O(INT0_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'h8B888BBBBBBBBBBB)) 
    INT0_carry_i_21
       (.I0(INT0_carry_i_28_n_0),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(ALU_DIN1[18]),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(ALU_DIN1[10]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry_i_21_n_0));
  LUT6 #(
    .INIT(64'h8B888BBBBBBBBBBB)) 
    INT0_carry_i_22
       (.I0(INT0_carry_i_17_n_0),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(ALU_DIN1[16]),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(ALU_DIN1[8]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry_i_22_n_0));
  LUT6 #(
    .INIT(64'h8B888BBBBBBBBBBB)) 
    INT0_carry_i_23
       (.I0(INT0_carry__0_i_17_n_0),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(ALU_DIN1[19]),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(ALU_DIN1[11]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry_i_23_n_0));
  LUT6 #(
    .INIT(64'h8B888BBBBBBBBBBB)) 
    INT0_carry_i_24
       (.I0(INT0_carry_i_20_n_0),
        .I1(INT0_carry__0_i_18_n_0),
        .I2(ALU_DIN1[17]),
        .I3(INT0_carry__2_i_13_n_0),
        .I4(ALU_DIN1[9]),
        .I5(INT0_carry__2_i_12_n_0),
        .O(INT0_carry_i_24_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry_i_25
       (.I0(INT0_carry_i_24_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry_i_18_n_0),
        .O(INT0_carry_i_25_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry_i_26
       (.I0(INT0_carry_i_22_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry_i_15_n_0),
        .O(INT0_carry_i_26_n_0));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    INT0_carry_i_27
       (.I0(ALU_DIN1[10]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[2]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[18]),
        .O(INT0_carry_i_27_n_0));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    INT0_carry_i_28
       (.I0(ALU_DIN1[14]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[6]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[22]),
        .O(INT0_carry_i_28_n_0));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    INT0_carry_i_29
       (.I0(ALU_DIN1[11]),
        .I1(INT0_carry__2_i_13_n_0),
        .I2(ALU_DIN1[3]),
        .I3(INT0_carry__2_i_12_n_0),
        .I4(ALU_DIN1[19]),
        .O(INT0_carry_i_29_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry_i_3
       (.I0(INT0_carry_i_11_n_0),
        .O(\custom_alu/fp2int/p_0_in [3]));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry_i_4
       (.I0(INT0_carry_i_12_n_0),
        .O(\custom_alu/fp2int/p_0_in [2]));
  LUT1 #(
    .INIT(2'h1)) 
    INT0_carry_i_5
       (.I0(INT0_carry_i_13_n_0),
        .O(\custom_alu/fp2int/p_0_in [1]));
  LUT6 #(
    .INIT(64'hFE7FFEFEFE7F7F7F)) 
    INT0_carry_i_6
       (.I0(INT0_carry_i_14_n_0),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[28]),
        .I3(ID_EX_Q[156]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I5(EX_RF_RD1[30]),
        .O(INT0_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'hBE82BEBEBE828282)) 
    INT0_carry_i_7
       (.I0(INT0_carry_i_15_n_0),
        .I1(ALU_DIN1[23]),
        .I2(ALU_DIN1[24]),
        .I3(INT0_carry_i_16_n_0),
        .I4(ALU_DIN1[25]),
        .I5(INT0_carry_i_17_n_0),
        .O(INT0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hBE82BEBEBE828282)) 
    INT0_carry_i_8
       (.I0(INT0_carry_i_18_n_0),
        .I1(ALU_DIN1[23]),
        .I2(ALU_DIN1[24]),
        .I3(INT0_carry_i_19_n_0),
        .I4(ALU_DIN1[25]),
        .I5(INT0_carry_i_20_n_0),
        .O(INT0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'hBBBEEEBE88822282)) 
    INT0_carry_i_9
       (.I0(INT0_carry_i_21_n_0),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD1[24]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(ID_EX_Q[150]),
        .I5(INT0_carry_i_22_n_0),
        .O(INT0_carry_i_9_n_0));
  OBUF \I_MEM_ADDR_OBUF[0]_inst 
       (.I(I_MEM_ADDR_OBUF[0]),
        .O(I_MEM_ADDR[0]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[0]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[0]),
        .I2(STALL_EN),
        .I3(IF_PC2[0]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[0] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[0]));
  OBUF \I_MEM_ADDR_OBUF[10]_inst 
       (.I(I_MEM_ADDR_OBUF[10]),
        .O(I_MEM_ADDR[10]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[10]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[10]),
        .I2(STALL_EN),
        .I3(IF_PC2[10]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[10] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[10]));
  OBUF \I_MEM_ADDR_OBUF[11]_inst 
       (.I(I_MEM_ADDR_OBUF[11]),
        .O(I_MEM_ADDR[11]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[11]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[11]),
        .I2(STALL_EN),
        .I3(IF_PC2[11]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[11] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[11]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[11]_inst_i_2 
       (.CI(\I_MEM_ADDR_OBUF[7]_inst_i_2_n_0 ),
        .CO({\I_MEM_ADDR_OBUF[11]_inst_i_2_n_0 ,\I_MEM_ADDR_OBUF[11]_inst_i_2_n_1 ,\I_MEM_ADDR_OBUF[11]_inst_i_2_n_2 ,\I_MEM_ADDR_OBUF[11]_inst_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ID_EX_Q[90:87]),
        .O(IF_PC2[11:8]),
        .S({\I_MEM_ADDR_OBUF[11]_inst_i_3_n_0 ,\I_MEM_ADDR_OBUF[11]_inst_i_4_n_0 ,\I_MEM_ADDR_OBUF[11]_inst_i_5_n_0 ,\I_MEM_ADDR_OBUF[11]_inst_i_6_n_0 }));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[11]_inst_i_3 
       (.I0(ID_EX_Q[90]),
        .I1(ID_EX_Q[137]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[11]),
        .O(\I_MEM_ADDR_OBUF[11]_inst_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[11]_inst_i_4 
       (.I0(ID_EX_Q[89]),
        .I1(ID_EX_Q[136]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[10]),
        .O(\I_MEM_ADDR_OBUF[11]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[11]_inst_i_5 
       (.I0(ID_EX_Q[88]),
        .I1(ID_EX_Q[135]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[9]),
        .O(\I_MEM_ADDR_OBUF[11]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[11]_inst_i_6 
       (.I0(ID_EX_Q[87]),
        .I1(ID_EX_Q[134]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[8]),
        .O(\I_MEM_ADDR_OBUF[11]_inst_i_6_n_0 ));
  OBUF \I_MEM_ADDR_OBUF[12]_inst 
       (.I(I_MEM_ADDR_OBUF[12]),
        .O(I_MEM_ADDR[12]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[12]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[12]),
        .I2(STALL_EN),
        .I3(IF_PC2[12]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[12] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[12]));
  OBUF \I_MEM_ADDR_OBUF[13]_inst 
       (.I(I_MEM_ADDR_OBUF[13]),
        .O(I_MEM_ADDR[13]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[13]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[13]),
        .I2(STALL_EN),
        .I3(IF_PC2[13]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[13] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[13]));
  OBUF \I_MEM_ADDR_OBUF[14]_inst 
       (.I(I_MEM_ADDR_OBUF[14]),
        .O(I_MEM_ADDR[14]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[14]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[14]),
        .I2(STALL_EN),
        .I3(IF_PC2[14]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[14] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[14]));
  OBUF \I_MEM_ADDR_OBUF[15]_inst 
       (.I(I_MEM_ADDR_OBUF[15]),
        .O(I_MEM_ADDR[15]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[15]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[15]),
        .I2(STALL_EN),
        .I3(IF_PC2[15]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[15] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[15]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[15]_inst_i_2 
       (.CI(\I_MEM_ADDR_OBUF[11]_inst_i_2_n_0 ),
        .CO({\I_MEM_ADDR_OBUF[15]_inst_i_2_n_0 ,\I_MEM_ADDR_OBUF[15]_inst_i_2_n_1 ,\I_MEM_ADDR_OBUF[15]_inst_i_2_n_2 ,\I_MEM_ADDR_OBUF[15]_inst_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ID_EX_Q[94:91]),
        .O(IF_PC2[15:12]),
        .S({\I_MEM_ADDR_OBUF[15]_inst_i_3_n_0 ,\I_MEM_ADDR_OBUF[15]_inst_i_4_n_0 ,\I_MEM_ADDR_OBUF[15]_inst_i_5_n_0 ,\I_MEM_ADDR_OBUF[15]_inst_i_6_n_0 }));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[15]_inst_i_3 
       (.I0(ID_EX_Q[94]),
        .I1(ID_EX_Q[141]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[15]),
        .O(\I_MEM_ADDR_OBUF[15]_inst_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[15]_inst_i_4 
       (.I0(ID_EX_Q[93]),
        .I1(ID_EX_Q[140]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[14]),
        .O(\I_MEM_ADDR_OBUF[15]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[15]_inst_i_5 
       (.I0(ID_EX_Q[92]),
        .I1(ID_EX_Q[139]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[13]),
        .O(\I_MEM_ADDR_OBUF[15]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[15]_inst_i_6 
       (.I0(ID_EX_Q[91]),
        .I1(ID_EX_Q[138]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[12]),
        .O(\I_MEM_ADDR_OBUF[15]_inst_i_6_n_0 ));
  OBUF \I_MEM_ADDR_OBUF[16]_inst 
       (.I(I_MEM_ADDR_OBUF[16]),
        .O(I_MEM_ADDR[16]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[16]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[16]),
        .I2(STALL_EN),
        .I3(IF_PC2[16]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[16] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[16]));
  OBUF \I_MEM_ADDR_OBUF[17]_inst 
       (.I(I_MEM_ADDR_OBUF[17]),
        .O(I_MEM_ADDR[17]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[17]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[17]),
        .I2(STALL_EN),
        .I3(IF_PC2[17]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[17] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[17]));
  OBUF \I_MEM_ADDR_OBUF[18]_inst 
       (.I(I_MEM_ADDR_OBUF[18]),
        .O(I_MEM_ADDR[18]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[18]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[18]),
        .I2(STALL_EN),
        .I3(IF_PC2[18]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[18] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[18]));
  OBUF \I_MEM_ADDR_OBUF[19]_inst 
       (.I(I_MEM_ADDR_OBUF[19]),
        .O(I_MEM_ADDR[19]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[19]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[19]),
        .I2(STALL_EN),
        .I3(IF_PC2[19]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[19] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[19]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[19]_inst_i_2 
       (.CI(\I_MEM_ADDR_OBUF[15]_inst_i_2_n_0 ),
        .CO({\I_MEM_ADDR_OBUF[19]_inst_i_2_n_0 ,\I_MEM_ADDR_OBUF[19]_inst_i_2_n_1 ,\I_MEM_ADDR_OBUF[19]_inst_i_2_n_2 ,\I_MEM_ADDR_OBUF[19]_inst_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ID_EX_Q[98:95]),
        .O(IF_PC2[19:16]),
        .S({\I_MEM_ADDR_OBUF[19]_inst_i_3_n_0 ,\I_MEM_ADDR_OBUF[19]_inst_i_4_n_0 ,\I_MEM_ADDR_OBUF[19]_inst_i_5_n_0 ,\I_MEM_ADDR_OBUF[19]_inst_i_6_n_0 }));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[19]_inst_i_3 
       (.I0(ID_EX_Q[98]),
        .I1(ID_EX_Q[145]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[19]),
        .O(\I_MEM_ADDR_OBUF[19]_inst_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[19]_inst_i_4 
       (.I0(ID_EX_Q[97]),
        .I1(ID_EX_Q[144]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[18]),
        .O(\I_MEM_ADDR_OBUF[19]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[19]_inst_i_5 
       (.I0(ID_EX_Q[96]),
        .I1(ID_EX_Q[143]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[17]),
        .O(\I_MEM_ADDR_OBUF[19]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[19]_inst_i_6 
       (.I0(ID_EX_Q[95]),
        .I1(ID_EX_Q[142]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[16]),
        .O(\I_MEM_ADDR_OBUF[19]_inst_i_6_n_0 ));
  OBUF \I_MEM_ADDR_OBUF[1]_inst 
       (.I(I_MEM_ADDR_OBUF[1]),
        .O(I_MEM_ADDR[1]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[1]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[1]),
        .I2(STALL_EN),
        .I3(IF_PC2[1]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[1] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[1]));
  OBUF \I_MEM_ADDR_OBUF[20]_inst 
       (.I(I_MEM_ADDR_OBUF[20]),
        .O(I_MEM_ADDR[20]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[20]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[20]),
        .I2(STALL_EN),
        .I3(IF_PC2[20]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[20] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[20]));
  OBUF \I_MEM_ADDR_OBUF[21]_inst 
       (.I(I_MEM_ADDR_OBUF[21]),
        .O(I_MEM_ADDR[21]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[21]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[21]),
        .I2(STALL_EN),
        .I3(IF_PC2[21]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[21] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[21]));
  OBUF \I_MEM_ADDR_OBUF[22]_inst 
       (.I(I_MEM_ADDR_OBUF[22]),
        .O(I_MEM_ADDR[22]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[22]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[22]),
        .I2(STALL_EN),
        .I3(IF_PC2[22]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[22] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[22]));
  OBUF \I_MEM_ADDR_OBUF[23]_inst 
       (.I(I_MEM_ADDR_OBUF[23]),
        .O(I_MEM_ADDR[23]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[23]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[23]),
        .I2(STALL_EN),
        .I3(IF_PC2[23]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[23] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[23]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[23]_inst_i_2 
       (.CI(\I_MEM_ADDR_OBUF[19]_inst_i_2_n_0 ),
        .CO({\I_MEM_ADDR_OBUF[23]_inst_i_2_n_0 ,\I_MEM_ADDR_OBUF[23]_inst_i_2_n_1 ,\I_MEM_ADDR_OBUF[23]_inst_i_2_n_2 ,\I_MEM_ADDR_OBUF[23]_inst_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ID_EX_Q[102:99]),
        .O(IF_PC2[23:20]),
        .S({\I_MEM_ADDR_OBUF[23]_inst_i_3_n_0 ,\I_MEM_ADDR_OBUF[23]_inst_i_4_n_0 ,\I_MEM_ADDR_OBUF[23]_inst_i_5_n_0 ,\I_MEM_ADDR_OBUF[23]_inst_i_6_n_0 }));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[23]_inst_i_3 
       (.I0(ID_EX_Q[102]),
        .I1(ID_EX_Q[149]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[23]),
        .O(\I_MEM_ADDR_OBUF[23]_inst_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[23]_inst_i_4 
       (.I0(ID_EX_Q[101]),
        .I1(ID_EX_Q[148]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[22]),
        .O(\I_MEM_ADDR_OBUF[23]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[23]_inst_i_5 
       (.I0(ID_EX_Q[100]),
        .I1(ID_EX_Q[147]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[21]),
        .O(\I_MEM_ADDR_OBUF[23]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[23]_inst_i_6 
       (.I0(ID_EX_Q[99]),
        .I1(ID_EX_Q[146]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[20]),
        .O(\I_MEM_ADDR_OBUF[23]_inst_i_6_n_0 ));
  OBUF \I_MEM_ADDR_OBUF[24]_inst 
       (.I(I_MEM_ADDR_OBUF[24]),
        .O(I_MEM_ADDR[24]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[24]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[24]),
        .I2(STALL_EN),
        .I3(IF_PC2[24]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[24] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[24]));
  OBUF \I_MEM_ADDR_OBUF[25]_inst 
       (.I(I_MEM_ADDR_OBUF[25]),
        .O(I_MEM_ADDR[25]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[25]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[25]),
        .I2(STALL_EN),
        .I3(IF_PC2[25]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[25] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[25]));
  OBUF \I_MEM_ADDR_OBUF[26]_inst 
       (.I(I_MEM_ADDR_OBUF[26]),
        .O(I_MEM_ADDR[26]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[26]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[26]),
        .I2(STALL_EN),
        .I3(IF_PC2[26]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[26] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[26]));
  OBUF \I_MEM_ADDR_OBUF[27]_inst 
       (.I(I_MEM_ADDR_OBUF[27]),
        .O(I_MEM_ADDR[27]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[27]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[27]),
        .I2(STALL_EN),
        .I3(IF_PC2[27]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[27] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[27]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[27]_inst_i_2 
       (.CI(\I_MEM_ADDR_OBUF[23]_inst_i_2_n_0 ),
        .CO({\I_MEM_ADDR_OBUF[27]_inst_i_2_n_0 ,\I_MEM_ADDR_OBUF[27]_inst_i_2_n_1 ,\I_MEM_ADDR_OBUF[27]_inst_i_2_n_2 ,\I_MEM_ADDR_OBUF[27]_inst_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ID_EX_Q[106:103]),
        .O(IF_PC2[27:24]),
        .S({\I_MEM_ADDR_OBUF[27]_inst_i_3_n_0 ,\I_MEM_ADDR_OBUF[27]_inst_i_4_n_0 ,\I_MEM_ADDR_OBUF[27]_inst_i_5_n_0 ,\I_MEM_ADDR_OBUF[27]_inst_i_6_n_0 }));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[27]_inst_i_3 
       (.I0(ID_EX_Q[106]),
        .I1(ID_EX_Q[153]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[27]),
        .O(\I_MEM_ADDR_OBUF[27]_inst_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[27]_inst_i_4 
       (.I0(ID_EX_Q[105]),
        .I1(ID_EX_Q[152]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[26]),
        .O(\I_MEM_ADDR_OBUF[27]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[27]_inst_i_5 
       (.I0(ID_EX_Q[104]),
        .I1(ID_EX_Q[151]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[25]),
        .O(\I_MEM_ADDR_OBUF[27]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[27]_inst_i_6 
       (.I0(ID_EX_Q[103]),
        .I1(ID_EX_Q[150]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[24]),
        .O(\I_MEM_ADDR_OBUF[27]_inst_i_6_n_0 ));
  OBUF \I_MEM_ADDR_OBUF[28]_inst 
       (.I(I_MEM_ADDR_OBUF[28]),
        .O(I_MEM_ADDR[28]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[28]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[28]),
        .I2(STALL_EN),
        .I3(IF_PC2[28]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[28] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[28]));
  OBUF \I_MEM_ADDR_OBUF[29]_inst 
       (.I(I_MEM_ADDR_OBUF[29]),
        .O(I_MEM_ADDR[29]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[29]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[29]),
        .I2(STALL_EN),
        .I3(IF_PC2[29]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[29] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[29]));
  OBUF \I_MEM_ADDR_OBUF[2]_inst 
       (.I(I_MEM_ADDR_OBUF[2]),
        .O(I_MEM_ADDR[2]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[2]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[2]),
        .I2(STALL_EN),
        .I3(IF_PC2[2]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[2] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[2]));
  OBUF \I_MEM_ADDR_OBUF[30]_inst 
       (.I(I_MEM_ADDR_OBUF[30]),
        .O(I_MEM_ADDR[30]));
  LUT6 #(
    .INIT(64'hFFFF00FFE4FFE4FF)) 
    \I_MEM_ADDR_OBUF[30]_inst_i_1 
       (.I0(EX_BR_TAKEN),
        .I1(\FF_IF_ID_PCADD/Q_reg_n_0_[30] ),
        .I2(IF_PC2[30]),
        .I3(RSTn_IBUF),
        .I4(ID_PC[30]),
        .I5(STALL_EN),
        .O(I_MEM_ADDR_OBUF[30]));
  OBUF \I_MEM_ADDR_OBUF[31]_inst 
       (.I(I_MEM_ADDR_OBUF[31]),
        .O(I_MEM_ADDR[31]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[31]),
        .I2(STALL_EN),
        .I3(IF_PC2[31]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[31] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[31]));
  LUT3 #(
    .INIT(8'h01)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_10 
       (.I0(STALL_COUNTER_Q[8]),
        .I1(STALL_COUNTER_Q[7]),
        .I2(STALL_COUNTER_Q[6]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_11 
       (.I0(STALL_COUNTER_Q[5]),
        .I1(STALL_COUNTER_Q[4]),
        .I2(STALL_COUNTER_Q[3]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8700000000008700)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_12 
       (.I0(\Q[79]_i_3_n_0 ),
        .I1(\Q[112]_i_2_n_0 ),
        .I2(STALL_COUNTER_Q[0]),
        .I3(\Q[9]_i_14_n_0 ),
        .I4(STALL_COUNTER_Q[1]),
        .I5(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_2 
       (.I0(LU_HAZARD),
        .I1(\stall_generator/CUSTOM_STALL ),
        .O(STALL_EN));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[31]_inst_i_3 
       (.CI(\I_MEM_ADDR_OBUF[27]_inst_i_2_n_0 ),
        .CO({\I_MEM_ADDR_OBUF[31]_inst_i_3_n_1 ,\I_MEM_ADDR_OBUF[31]_inst_i_3_n_2 ,\I_MEM_ADDR_OBUF[31]_inst_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,ID_EX_Q[109:107]}),
        .O(IF_PC2[31:28]),
        .S({\I_MEM_ADDR_OBUF[31]_inst_i_5_n_0 ,\I_MEM_ADDR_OBUF[31]_inst_i_6_n_0 ,\I_MEM_ADDR_OBUF[31]_inst_i_7_n_0 ,\I_MEM_ADDR_OBUF[31]_inst_i_8_n_0 }));
  CARRY4 \I_MEM_ADDR_OBUF[31]_inst_i_4 
       (.CI(\<const0> ),
        .CO({\stall_generator/CUSTOM_STALL ,\I_MEM_ADDR_OBUF[31]_inst_i_4_n_1 ,\I_MEM_ADDR_OBUF[31]_inst_i_4_n_2 ,\I_MEM_ADDR_OBUF[31]_inst_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const1> ,\<const1> ,\<const1> ,\<const1> }),
        .S({\I_MEM_ADDR_OBUF[31]_inst_i_9_n_0 ,\I_MEM_ADDR_OBUF[31]_inst_i_10_n_0 ,\I_MEM_ADDR_OBUF[31]_inst_i_11_n_0 ,\I_MEM_ADDR_OBUF[31]_inst_i_12_n_0 }));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_5 
       (.I0(ID_EX_Q[110]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[31]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_6 
       (.I0(ID_EX_Q[109]),
        .I1(ID_EX_Q[156]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[30]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_7 
       (.I0(ID_EX_Q[108]),
        .I1(ID_EX_Q[155]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[29]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_8 
       (.I0(ID_EX_Q[107]),
        .I1(ID_EX_Q[154]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[28]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_8_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \I_MEM_ADDR_OBUF[31]_inst_i_9 
       (.I0(STALL_COUNTER_Q[9]),
        .O(\I_MEM_ADDR_OBUF[31]_inst_i_9_n_0 ));
  OBUF \I_MEM_ADDR_OBUF[3]_inst 
       (.I(I_MEM_ADDR_OBUF[3]),
        .O(I_MEM_ADDR[3]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[3]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[3]),
        .I2(STALL_EN),
        .I3(IF_PC2[3]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[3] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[3]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[3]_inst_i_2 
       (.CI(\<const0> ),
        .CO({\I_MEM_ADDR_OBUF[3]_inst_i_2_n_0 ,\I_MEM_ADDR_OBUF[3]_inst_i_2_n_1 ,\I_MEM_ADDR_OBUF[3]_inst_i_2_n_2 ,\I_MEM_ADDR_OBUF[3]_inst_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({ID_EX_Q[82:80],\<const0> }),
        .O(IF_PC2[3:0]),
        .S({\I_MEM_ADDR_OBUF[3]_inst_i_3_n_0 ,\I_MEM_ADDR_OBUF[3]_inst_i_4_n_0 ,\I_MEM_ADDR_OBUF[3]_inst_i_5_n_0 ,p_0_in}));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[3]_inst_i_3 
       (.I0(ID_EX_Q[82]),
        .I1(ID_EX_Q[129]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[3]),
        .O(\I_MEM_ADDR_OBUF[3]_inst_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[3]_inst_i_4 
       (.I0(ID_EX_Q[81]),
        .I1(ID_EX_Q[128]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[2]),
        .O(\I_MEM_ADDR_OBUF[3]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[3]_inst_i_5 
       (.I0(ID_EX_Q[80]),
        .I1(ID_EX_Q[127]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[1]),
        .O(\I_MEM_ADDR_OBUF[3]_inst_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \I_MEM_ADDR_OBUF[3]_inst_i_6 
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I2(ID_EX_Q[126]),
        .O(p_0_in));
  OBUF \I_MEM_ADDR_OBUF[4]_inst 
       (.I(I_MEM_ADDR_OBUF[4]),
        .O(I_MEM_ADDR[4]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[4]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[4]),
        .I2(STALL_EN),
        .I3(IF_PC2[4]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[4] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[4]));
  OBUF \I_MEM_ADDR_OBUF[5]_inst 
       (.I(I_MEM_ADDR_OBUF[5]),
        .O(I_MEM_ADDR[5]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[5]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[5]),
        .I2(STALL_EN),
        .I3(IF_PC2[5]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[5] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[5]));
  OBUF \I_MEM_ADDR_OBUF[6]_inst 
       (.I(I_MEM_ADDR_OBUF[6]),
        .O(I_MEM_ADDR[6]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[6]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[6]),
        .I2(STALL_EN),
        .I3(IF_PC2[6]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[6] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[6]));
  OBUF \I_MEM_ADDR_OBUF[7]_inst 
       (.I(I_MEM_ADDR_OBUF[7]),
        .O(I_MEM_ADDR[7]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[7]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[7]),
        .I2(STALL_EN),
        .I3(IF_PC2[7]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[7] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[7]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \I_MEM_ADDR_OBUF[7]_inst_i_2 
       (.CI(\I_MEM_ADDR_OBUF[3]_inst_i_2_n_0 ),
        .CO({\I_MEM_ADDR_OBUF[7]_inst_i_2_n_0 ,\I_MEM_ADDR_OBUF[7]_inst_i_2_n_1 ,\I_MEM_ADDR_OBUF[7]_inst_i_2_n_2 ,\I_MEM_ADDR_OBUF[7]_inst_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(ID_EX_Q[86:83]),
        .O(IF_PC2[7:4]),
        .S({\I_MEM_ADDR_OBUF[7]_inst_i_3_n_0 ,\I_MEM_ADDR_OBUF[7]_inst_i_4_n_0 ,\I_MEM_ADDR_OBUF[7]_inst_i_5_n_0 ,\I_MEM_ADDR_OBUF[7]_inst_i_6_n_0 }));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[7]_inst_i_3 
       (.I0(ID_EX_Q[86]),
        .I1(ID_EX_Q[133]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[7]),
        .O(\I_MEM_ADDR_OBUF[7]_inst_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[7]_inst_i_4 
       (.I0(ID_EX_Q[85]),
        .I1(ID_EX_Q[132]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[6]),
        .O(\I_MEM_ADDR_OBUF[7]_inst_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[7]_inst_i_5 
       (.I0(ID_EX_Q[84]),
        .I1(ID_EX_Q[131]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[5]),
        .O(\I_MEM_ADDR_OBUF[7]_inst_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56A6)) 
    \I_MEM_ADDR_OBUF[7]_inst_i_6 
       (.I0(ID_EX_Q[83]),
        .I1(ID_EX_Q[130]),
        .I2(\FF_JALR_EN/Q_reg_n_0_[0] ),
        .I3(EX_RF_RD1[4]),
        .O(\I_MEM_ADDR_OBUF[7]_inst_i_6_n_0 ));
  OBUF \I_MEM_ADDR_OBUF[8]_inst 
       (.I(I_MEM_ADDR_OBUF[8]),
        .O(I_MEM_ADDR[8]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[8]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[8]),
        .I2(STALL_EN),
        .I3(IF_PC2[8]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[8] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[8]));
  OBUF \I_MEM_ADDR_OBUF[9]_inst 
       (.I(I_MEM_ADDR_OBUF[9]),
        .O(I_MEM_ADDR[9]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \I_MEM_ADDR_OBUF[9]_inst_i_1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[9]),
        .I2(STALL_EN),
        .I3(IF_PC2[9]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[9] ),
        .I5(EX_BR_TAKEN),
        .O(I_MEM_ADDR_OBUF[9]));
  OBUF I_MEM_CSN_OBUF_inst
       (.I(\<const0> ),
        .O(I_MEM_CSN));
  IBUF \I_MEM_DOUT_IBUF[10]_inst 
       (.I(I_MEM_DOUT[10]),
        .O(I_MEM_DOUT_IBUF[10]));
  IBUF \I_MEM_DOUT_IBUF[11]_inst 
       (.I(I_MEM_DOUT[11]),
        .O(I_MEM_DOUT_IBUF[11]));
  IBUF \I_MEM_DOUT_IBUF[12]_inst 
       (.I(I_MEM_DOUT[12]),
        .O(I_MEM_DOUT_IBUF[12]));
  IBUF \I_MEM_DOUT_IBUF[13]_inst 
       (.I(I_MEM_DOUT[13]),
        .O(I_MEM_DOUT_IBUF[13]));
  IBUF \I_MEM_DOUT_IBUF[14]_inst 
       (.I(I_MEM_DOUT[14]),
        .O(I_MEM_DOUT_IBUF[14]));
  IBUF \I_MEM_DOUT_IBUF[15]_inst 
       (.I(I_MEM_DOUT[15]),
        .O(CRF_RA1_OBUF[0]));
  IBUF \I_MEM_DOUT_IBUF[16]_inst 
       (.I(I_MEM_DOUT[16]),
        .O(CRF_RA1_OBUF[1]));
  IBUF \I_MEM_DOUT_IBUF[17]_inst 
       (.I(I_MEM_DOUT[17]),
        .O(CRF_RA1_OBUF[2]));
  IBUF \I_MEM_DOUT_IBUF[18]_inst 
       (.I(I_MEM_DOUT[18]),
        .O(CRF_RA1_OBUF[3]));
  IBUF \I_MEM_DOUT_IBUF[19]_inst 
       (.I(I_MEM_DOUT[19]),
        .O(CRF_RA1_OBUF[4]));
  IBUF \I_MEM_DOUT_IBUF[20]_inst 
       (.I(I_MEM_DOUT[20]),
        .O(CRF_RA2_OBUF[0]));
  IBUF \I_MEM_DOUT_IBUF[21]_inst 
       (.I(I_MEM_DOUT[21]),
        .O(CRF_RA2_OBUF[1]));
  IBUF \I_MEM_DOUT_IBUF[22]_inst 
       (.I(I_MEM_DOUT[22]),
        .O(CRF_RA2_OBUF[2]));
  IBUF \I_MEM_DOUT_IBUF[23]_inst 
       (.I(I_MEM_DOUT[23]),
        .O(CRF_RA2_OBUF[3]));
  IBUF \I_MEM_DOUT_IBUF[24]_inst 
       (.I(I_MEM_DOUT[24]),
        .O(CRF_RA2_OBUF[4]));
  IBUF \I_MEM_DOUT_IBUF[25]_inst 
       (.I(I_MEM_DOUT[25]),
        .O(I_MEM_DOUT_IBUF[25]));
  IBUF \I_MEM_DOUT_IBUF[26]_inst 
       (.I(I_MEM_DOUT[26]),
        .O(I_MEM_DOUT_IBUF[26]));
  IBUF \I_MEM_DOUT_IBUF[27]_inst 
       (.I(I_MEM_DOUT[27]),
        .O(I_MEM_DOUT_IBUF[27]));
  IBUF \I_MEM_DOUT_IBUF[28]_inst 
       (.I(I_MEM_DOUT[28]),
        .O(I_MEM_DOUT_IBUF[28]));
  IBUF \I_MEM_DOUT_IBUF[29]_inst 
       (.I(I_MEM_DOUT[29]),
        .O(I_MEM_DOUT_IBUF[29]));
  IBUF \I_MEM_DOUT_IBUF[2]_inst 
       (.I(I_MEM_DOUT[2]),
        .O(I_MEM_DOUT_IBUF[2]));
  IBUF \I_MEM_DOUT_IBUF[30]_inst 
       (.I(I_MEM_DOUT[30]),
        .O(I_MEM_DOUT_IBUF[30]));
  IBUF \I_MEM_DOUT_IBUF[31]_inst 
       (.I(I_MEM_DOUT[31]),
        .O(I_MEM_DOUT_IBUF[31]));
  IBUF \I_MEM_DOUT_IBUF[3]_inst 
       (.I(I_MEM_DOUT[3]),
        .O(I_MEM_DOUT_IBUF[3]));
  IBUF \I_MEM_DOUT_IBUF[4]_inst 
       (.I(I_MEM_DOUT[4]),
        .O(I_MEM_DOUT_IBUF[4]));
  IBUF \I_MEM_DOUT_IBUF[5]_inst 
       (.I(I_MEM_DOUT[5]),
        .O(I_MEM_DOUT_IBUF[5]));
  IBUF \I_MEM_DOUT_IBUF[6]_inst 
       (.I(I_MEM_DOUT[6]),
        .O(I_MEM_DOUT_IBUF[6]));
  IBUF \I_MEM_DOUT_IBUF[7]_inst 
       (.I(I_MEM_DOUT[7]),
        .O(I_MEM_DOUT_IBUF[7]));
  IBUF \I_MEM_DOUT_IBUF[8]_inst 
       (.I(I_MEM_DOUT[8]),
        .O(I_MEM_DOUT_IBUF[8]));
  IBUF \I_MEM_DOUT_IBUF[9]_inst 
       (.I(I_MEM_DOUT[9]),
        .O(I_MEM_DOUT_IBUF[9]));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_1
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[22]),
        .O(PSUM0__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry__0_i_10
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM0__0_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry__0_i_10__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM0__0_carry__0_i_10__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry__0_i_10__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(ALU_DIN2[2]),
        .O(PSUM0__0_carry__0_i_10__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry__0_i_10__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(ALU_DIN2[2]),
        .O(PSUM0__0_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry__0_i_11
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[17]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[96]),
        .O(PSUM0__0_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry__0_i_11__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[17]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[96]),
        .O(PSUM0__0_carry__0_i_11__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry__0_i_11__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(ALU_DIN2[1]),
        .O(PSUM0__0_carry__0_i_11__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry__0_i_11__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(ALU_DIN2[1]),
        .O(PSUM0__0_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry__0_i_12
       (.I0(EX_RF_RD1[2]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[128]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM0__0_carry__0_i_12_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry__0_i_12__0
       (.I0(EX_RF_RD1[18]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[144]),
        .I3(ALU_DIN2[2]),
        .O(PSUM0__0_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM0__0_carry__0_i_12__1
       (.I0(ID_EX_Q[144]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[18]),
        .I3(ID_EX_Q[97]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[18]),
        .O(PSUM0__0_carry__0_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h47FF)) 
    PSUM0__0_carry__0_i_12__2
       (.I0(ID_EX_Q[128]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[2]),
        .I3(ALU_DIN2[2]),
        .O(PSUM0__0_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_1__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[6]),
        .O(PSUM0__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_1__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[22]),
        .O(PSUM0__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_1__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[6]),
        .O(PSUM0__0_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_2
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[21]),
        .O(PSUM0__0_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_2__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[5]),
        .O(PSUM0__0_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_2__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[21]),
        .O(PSUM0__0_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_2__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[5]),
        .O(PSUM0__0_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_3
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[20]),
        .O(PSUM0__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_3__0
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[4]),
        .O(PSUM0__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_3__1
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[4]),
        .O(PSUM0__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_3__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[20]),
        .O(PSUM0__0_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_4
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[19]),
        .O(PSUM0__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_4__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[3]),
        .O(PSUM0__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_4__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[19]),
        .O(PSUM0__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__0_i_4__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[3]),
        .O(PSUM0__0_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_5
       (.I0(PSUM0__0_carry__0_i_1_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM0__0_carry__0_i_9_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_5__0
       (.I0(PSUM0__0_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM0__0_carry__0_i_9__0_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_5__1
       (.I0(PSUM0__0_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM0__0_carry__0_i_9__1_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_5__2
       (.I0(PSUM0__0_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM0__0_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_6
       (.I0(PSUM0__0_carry__0_i_2_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM0__0_carry__0_i_10_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_6__0
       (.I0(PSUM0__0_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM0__0_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_6__1
       (.I0(PSUM0__0_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM0__0_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_6__2
       (.I0(PSUM0__0_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM0__0_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM0__0_carry__0_i_7
       (.I0(PSUM0__0_carry__0_i_3_n_0),
        .I1(PSUM0__0_carry__0_i_11_n_0),
        .I2(ALU_DIN2[18]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM0__0_carry__0_i_7__0
       (.I0(PSUM0__0_carry__0_i_3__0_n_0),
        .I1(PSUM0__0_carry__0_i_11__2_n_0),
        .I2(ALU_DIN2[2]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM0__0_carry__0_i_7__1
       (.I0(PSUM0__0_carry__0_i_3__1_n_0),
        .I1(PSUM0__0_carry__0_i_11__0_n_0),
        .I2(ALU_DIN2[18]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM0__0_carry__0_i_7__2
       (.I0(PSUM0__0_carry__0_i_3__2_n_0),
        .I1(PSUM0__0_carry__0_i_11__1_n_0),
        .I2(ALU_DIN2[2]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_8
       (.I0(PSUM0__0_carry__0_i_4_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[19]),
        .I3(PSUM0__0_carry__0_i_12__1_n_0),
        .I4(ALU_DIN1[20]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_8__0
       (.I0(PSUM0__0_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[3]),
        .I3(PSUM0__0_carry__0_i_12__2_n_0),
        .I4(ALU_DIN1[4]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_8__1
       (.I0(PSUM0__0_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[3]),
        .I3(PSUM0__0_carry__0_i_12_n_0),
        .I4(ALU_DIN1[4]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__0_carry__0_i_8__2
       (.I0(PSUM0__0_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[19]),
        .I3(PSUM0__0_carry__0_i_12__0_n_0),
        .I4(ALU_DIN1[20]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry__0_i_9
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM0__0_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry__0_i_9__0
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM0__0_carry__0_i_9__0_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry__0_i_9__1
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(ALU_DIN2[2]),
        .O(PSUM0__0_carry__0_i_9__1_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry__0_i_9__2
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(ALU_DIN2[2]),
        .O(PSUM0__0_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM0__0_carry__1_i_1
       (.I0(ID_EX_Q[97]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[18]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[17]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__0_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM0__0_carry__1_i_1__0
       (.I0(ID_EX_Q[97]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[18]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[17]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__0_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM0__0_carry__1_i_1__1
       (.I0(ALU_DIN2[2]),
        .I1(ID_EX_Q[148]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[22]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__0_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM0__0_carry__1_i_1__2
       (.I0(ALU_DIN2[2]),
        .I1(ID_EX_Q[132]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[6]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__0_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__1_i_2
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__0_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__1_i_2__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__0_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__1_i_2__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__0_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__0_carry__1_i_2__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__0_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM0__0_carry__1_i_3
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[96]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[18]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__0_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM0__0_carry__1_i_3__0
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[96]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[18]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__0_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM0__0_carry__1_i_3__1
       (.I0(ALU_DIN2[1]),
        .I1(EX_RF_RD1[22]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[148]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__0_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM0__0_carry__1_i_3__2
       (.I0(ALU_DIN2[1]),
        .I1(EX_RF_RD1[6]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[132]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__0_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__0_carry__1_i_4
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[18]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[17]),
        .O(PSUM0__0_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__0_carry__1_i_4__0
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[18]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[17]),
        .O(PSUM0__0_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__0_carry__1_i_4__1
       (.I0(ALU_DIN2[0]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[2]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[1]),
        .O(PSUM0__0_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__0_carry__1_i_4__2
       (.I0(ALU_DIN2[0]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[2]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[1]),
        .O(PSUM0__0_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_1
       (.I0(ALU_DIN2[17]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[18]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_1__0
       (.I0(ALU_DIN2[17]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[18]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[16]),
        .O(PSUM0__0_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_1__1
       (.I0(ALU_DIN2[1]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[2]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_1__2
       (.I0(ALU_DIN2[1]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[2]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[0]),
        .O(PSUM0__0_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h1DFFE200E200E200)) 
    PSUM0__0_carry_i_2
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[96]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[18]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__0_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h57F7A808A808A808)) 
    PSUM0__0_carry_i_2__0
       (.I0(ALU_DIN2[1]),
        .I1(EX_RF_RD1[1]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[127]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM0__0_carry_i_2__1
       (.I0(ID_EX_Q[96]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[17]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[18]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM0__0_carry_i_2__2
       (.I0(ALU_DIN2[1]),
        .I1(ID_EX_Q[143]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[17]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__0_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM0__0_carry_i_3
       (.I0(ID_EX_Q[95]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[16]),
        .I3(ID_EX_Q[143]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[17]),
        .O(PSUM0__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM0__0_carry_i_3__0
       (.I0(ID_EX_Q[95]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[16]),
        .I3(ID_EX_Q[127]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[1]),
        .O(PSUM0__0_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM0__0_carry_i_3__1
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[143]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[17]),
        .O(PSUM0__0_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM0__0_carry_i_3__2
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[127]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[1]),
        .O(PSUM0__0_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__0_carry_i_4
       (.I0(ALU_DIN1[18]),
        .I1(PSUM0__0_carry_i_8_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[18]),
        .O(PSUM0__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__0_carry_i_4__0
       (.I0(ALU_DIN1[2]),
        .I1(PSUM0__0_carry_i_8__2_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[2]),
        .O(PSUM0__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__0_carry_i_4__1
       (.I0(ALU_DIN1[2]),
        .I1(PSUM0__0_carry_i_8__0_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[18]),
        .O(PSUM0__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__0_carry_i_4__2
       (.I0(ALU_DIN1[18]),
        .I1(PSUM0__0_carry_i_8__1_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[2]),
        .O(PSUM0__0_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_5
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[18]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[18]),
        .O(PSUM0__0_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_5__0
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[2]),
        .O(PSUM0__0_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_5__1
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[18]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[2]),
        .O(PSUM0__0_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__0_carry_i_5__2
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[18]),
        .O(PSUM0__0_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM0__0_carry_i_6
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[17]),
        .I2(ID_EX_Q[96]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[17]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__0_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM0__0_carry_i_6__0
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[1]),
        .I2(ID_EX_Q[96]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[17]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__0_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM0__0_carry_i_6__1
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[143]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[17]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__0_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM0__0_carry_i_6__2
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[127]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[1]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__0_carry_i_6__2_n_0));
  LUT4 #(
    .INIT(16'hB800)) 
    PSUM0__0_carry_i_7
       (.I0(ID_EX_Q[126]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[0]),
        .I3(ALU_DIN2[0]),
        .O(PSUM0__0_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    PSUM0__0_carry_i_7__0
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(ALU_DIN2[0]),
        .O(PSUM0__0_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM0__0_carry_i_7__1
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM0__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM0__0_carry_i_7__2
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM0__0_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry_i_8
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM0__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__0_carry_i_8__0
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM0__0_carry_i_8__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry_i_8__1
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(ALU_DIN2[0]),
        .O(PSUM0__0_carry_i_8__1_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__0_carry_i_8__2
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(ALU_DIN2[0]),
        .O(PSUM0__0_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_1
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[22]),
        .O(PSUM0__30_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_10
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM0__30_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_10__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM0__30_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_10__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM0__30_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_10__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM0__30_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_11
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[20]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[99]),
        .O(PSUM0__30_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_11__0
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM0__30_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_11__1
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM0__30_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM0__30_carry__0_i_11__2
       (.I0(ID_EX_Q[146]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[20]),
        .I3(ID_EX_Q[99]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[20]),
        .O(PSUM0__30_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_12
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM0__30_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_12__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM0__30_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_12__1
       (.I0(EX_RF_RD1[18]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[144]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM0__30_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_12__2
       (.I0(EX_RF_RD1[2]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[128]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM0__30_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_1__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[6]),
        .O(PSUM0__30_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_1__1
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[22]),
        .O(PSUM0__30_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_1__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[6]),
        .O(PSUM0__30_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[5]),
        .O(PSUM0__30_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_2__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[21]),
        .O(PSUM0__30_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_2__1
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[5]),
        .O(PSUM0__30_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_2__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[21]),
        .O(PSUM0__30_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_3
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[20]),
        .O(PSUM0__30_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_3__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[4]),
        .O(PSUM0__30_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_3__1
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[20]),
        .O(PSUM0__30_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_3__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[4]),
        .O(PSUM0__30_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_4
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[19]),
        .O(PSUM0__30_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_4__0
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[3]),
        .O(PSUM0__30_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_4__1
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[3]),
        .O(PSUM0__30_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__0_i_4__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[19]),
        .O(PSUM0__30_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_5
       (.I0(PSUM0__30_carry__0_i_1_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM0__30_carry__0_i_9__1_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_5__0
       (.I0(PSUM0__30_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM0__30_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_5__1
       (.I0(PSUM0__30_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM0__30_carry__0_i_9_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_5__2
       (.I0(PSUM0__30_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM0__30_carry__0_i_9__0_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_6
       (.I0(PSUM0__30_carry__0_i_2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM0__30_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_6__0
       (.I0(PSUM0__30_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM0__30_carry__0_i_10_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_6__1
       (.I0(PSUM0__30_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM0__30_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_6__2
       (.I0(PSUM0__30_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM0__30_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_7
       (.I0(PSUM0__30_carry__0_i_3__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[4]),
        .I3(PSUM0__30_carry__0_i_11__1_n_0),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM0__30_carry__0_i_7__0
       (.I0(PSUM0__30_carry__0_i_3_n_0),
        .I1(PSUM0__30_carry__0_i_11__2_n_0),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM0__30_carry__0_i_7__1
       (.I0(PSUM0__30_carry__0_i_3__0_n_0),
        .I1(PSUM0__30_carry__0_i_11_n_0),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_7__2
       (.I0(PSUM0__30_carry__0_i_3__1_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[20]),
        .I3(PSUM0__30_carry__0_i_11__0_n_0),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A6A6A959595)) 
    PSUM0__30_carry__0_i_8
       (.I0(PSUM0__30_carry__0_i_4_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[19]),
        .I3(ALU_DIN2[21]),
        .I4(ALU_DIN1[18]),
        .I5(PSUM0__30_carry__0_i_12_n_0),
        .O(PSUM0__30_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_8__0
       (.I0(PSUM0__30_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[3]),
        .I3(PSUM0__30_carry__0_i_12__2_n_0),
        .I4(ALU_DIN1[4]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A6A6A959595)) 
    PSUM0__30_carry__0_i_8__1
       (.I0(PSUM0__30_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[3]),
        .I3(ALU_DIN2[21]),
        .I4(ALU_DIN1[2]),
        .I5(PSUM0__30_carry__0_i_12__0_n_0),
        .O(PSUM0__30_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM0__30_carry__0_i_8__2
       (.I0(PSUM0__30_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[19]),
        .I3(PSUM0__30_carry__0_i_12__1_n_0),
        .I4(ALU_DIN1[20]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_9
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM0__30_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry__0_i_9__0
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM0__30_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM0__30_carry__0_i_9__1
       (.I0(ID_EX_Q[147]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[21]),
        .I3(ID_EX_Q[100]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[21]),
        .O(PSUM0__30_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM0__30_carry__0_i_9__2
       (.I0(ID_EX_Q[131]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[5]),
        .I3(ID_EX_Q[84]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[5]),
        .O(PSUM0__30_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM0__30_carry__1_i_1
       (.I0(ID_EX_Q[100]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[21]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[20]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__30_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM0__30_carry__1_i_1__0
       (.I0(ID_EX_Q[100]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[21]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[20]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__30_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM0__30_carry__1_i_1__1
       (.I0(ALU_DIN2[5]),
        .I1(ID_EX_Q[148]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[22]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__30_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM0__30_carry__1_i_1__2
       (.I0(ALU_DIN2[5]),
        .I1(ID_EX_Q[132]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[6]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__30_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__1_i_2
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__30_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__1_i_2__0
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__30_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__1_i_2__1
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__30_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM0__30_carry__1_i_2__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__30_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM0__30_carry__1_i_3
       (.I0(EX_RF_RD2[20]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[99]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[21]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__30_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM0__30_carry__1_i_3__0
       (.I0(EX_RF_RD2[20]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[99]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[21]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__30_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM0__30_carry__1_i_3__1
       (.I0(ALU_DIN2[4]),
        .I1(EX_RF_RD1[22]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[148]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[23]),
        .O(PSUM0__30_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM0__30_carry__1_i_3__2
       (.I0(ALU_DIN2[4]),
        .I1(EX_RF_RD1[6]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[132]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[7]),
        .O(PSUM0__30_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__30_carry__1_i_4
       (.I0(ALU_DIN2[19]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[21]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[20]),
        .O(PSUM0__30_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__30_carry__1_i_4__0
       (.I0(ALU_DIN2[3]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[4]),
        .O(PSUM0__30_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__30_carry__1_i_4__1
       (.I0(ALU_DIN2[19]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[21]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[20]),
        .O(PSUM0__30_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM0__30_carry__1_i_4__2
       (.I0(ALU_DIN2[3]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[4]),
        .O(PSUM0__30_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_1
       (.I0(ALU_DIN2[20]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_1__0
       (.I0(ALU_DIN2[4]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_1__1
       (.I0(ALU_DIN2[20]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[19]),
        .O(PSUM0__30_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_1__2
       (.I0(ALU_DIN2[4]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[3]),
        .O(PSUM0__30_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM0__30_carry_i_2
       (.I0(ID_EX_Q[99]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[20]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[21]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__30_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM0__30_carry_i_2__0
       (.I0(ID_EX_Q[99]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[20]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[21]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__30_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM0__30_carry_i_2__1
       (.I0(ALU_DIN2[4]),
        .I1(ID_EX_Q[143]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[17]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__30_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM0__30_carry_i_2__2
       (.I0(ALU_DIN2[4]),
        .I1(ID_EX_Q[127]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[1]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__30_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM0__30_carry_i_3
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ID_EX_Q[143]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[17]),
        .O(PSUM0__30_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM0__30_carry_i_3__0
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ID_EX_Q[127]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[1]),
        .O(PSUM0__30_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM0__30_carry_i_3__1
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[143]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[17]),
        .O(PSUM0__30_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM0__30_carry_i_3__2
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[127]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[1]),
        .O(PSUM0__30_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__30_carry_i_4
       (.I0(ALU_DIN1[18]),
        .I1(PSUM0__30_carry_i_8__1_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[21]),
        .O(PSUM0__30_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__30_carry_i_4__0
       (.I0(ALU_DIN1[2]),
        .I1(PSUM0__30_carry_i_8__2_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[5]),
        .O(PSUM0__30_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__30_carry_i_4__1
       (.I0(ALU_DIN1[2]),
        .I1(PSUM0__30_carry_i_8_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[21]),
        .O(PSUM0__30_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM0__30_carry_i_4__2
       (.I0(ALU_DIN1[18]),
        .I1(PSUM0__30_carry_i_8__0_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[5]),
        .O(PSUM0__30_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_5
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[21]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[18]),
        .O(PSUM0__30_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_5__0
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[21]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[2]),
        .O(PSUM0__30_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_5__1
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[5]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[18]),
        .O(PSUM0__30_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM0__30_carry_i_5__2
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[5]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[2]),
        .O(PSUM0__30_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM0__30_carry_i_6
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[20]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__30_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM0__30_carry_i_6__0
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[20]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__30_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM0__30_carry_i_6__1
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[143]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[17]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__30_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM0__30_carry_i_6__2
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[127]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[1]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__30_carry_i_6__2_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    PSUM0__30_carry_i_7
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(ALU_DIN2[3]),
        .O(PSUM0__30_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM0__30_carry_i_7__0
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM0__30_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    PSUM0__30_carry_i_7__1
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(ALU_DIN2[3]),
        .O(PSUM0__30_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM0__30_carry_i_7__2
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM0__30_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__30_carry_i_8
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM0__30_carry_i_8_n_0));
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM0__30_carry_i_8__0
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(ALU_DIN2[3]),
        .O(PSUM0__30_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM0__30_carry_i_8__1
       (.I0(ID_EX_Q[145]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[19]),
        .I3(ID_EX_Q[98]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[19]),
        .O(PSUM0__30_carry_i_8__1_n_0));
  LUT4 #(
    .INIT(16'h47FF)) 
    PSUM0__30_carry_i_8__2
       (.I0(ID_EX_Q[129]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[3]),
        .I3(ALU_DIN2[3]),
        .O(PSUM0__30_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__0_i_1
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM0__60_carry__0_i_9_n_0),
        .I5(PSUM0__60_carry__0_i_10_n_0),
        .O(PSUM0__60_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_10
       (.I0(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_7 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[17]),
        .O(PSUM0__60_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_10__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_7 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[1]),
        .O(PSUM0__60_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_10__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_7 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[17]),
        .O(PSUM0__60_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_10__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_7 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[1]),
        .O(PSUM0__60_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_11
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_7 ),
        .O(PSUM0__60_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_11__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_7 ),
        .O(PSUM0__60_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_11__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_7 ),
        .O(PSUM0__60_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_11__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_7 ),
        .O(PSUM0__60_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_12
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[19]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_1 ),
        .O(PSUM0__60_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_12__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[3]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_1 ),
        .O(PSUM0__60_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_12__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[19]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_1 ),
        .O(PSUM0__60_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_12__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[3]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_1 ),
        .O(PSUM0__60_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_13
       (.I0(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_6 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[18]),
        .O(PSUM0__60_carry__0_i_13_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_13__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_6 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[2]),
        .O(PSUM0__60_carry__0_i_13__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_13__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_6 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[18]),
        .O(PSUM0__60_carry__0_i_13__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__0_i_13__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_6 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[2]),
        .O(PSUM0__60_carry__0_i_13__2_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM0__60_carry__0_i_14
       (.I0(ALU_DIN1[17]),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[22]),
        .I5(PSUM0__60_carry__0_i_11_n_0),
        .O(PSUM0__60_carry__0_i_14_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM0__60_carry__0_i_14__0
       (.I0(ALU_DIN1[1]),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[22]),
        .I5(PSUM0__60_carry__0_i_11__0_n_0),
        .O(PSUM0__60_carry__0_i_14__0_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM0__60_carry__0_i_14__1
       (.I0(ALU_DIN1[17]),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[6]),
        .I5(PSUM0__60_carry__0_i_11__1_n_0),
        .O(PSUM0__60_carry__0_i_14__1_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM0__60_carry__0_i_14__2
       (.I0(ALU_DIN1[1]),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[6]),
        .I5(PSUM0__60_carry__0_i_11__2_n_0),
        .O(PSUM0__60_carry__0_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_15
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[16]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_4 ),
        .O(PSUM0__60_carry__0_i_15_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_15__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[0]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_4 ),
        .O(PSUM0__60_carry__0_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_15__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[16]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_4 ),
        .O(PSUM0__60_carry__0_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_15__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[0]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_4 ),
        .O(PSUM0__60_carry__0_i_15__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__0_i_1__0
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM0__60_carry__0_i_9__0_n_0),
        .I5(PSUM0__60_carry__0_i_10__0_n_0),
        .O(PSUM0__60_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__0_i_1__1
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM0__60_carry__0_i_9__1_n_0),
        .I5(PSUM0__60_carry__0_i_10__1_n_0),
        .O(PSUM0__60_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__0_i_1__2
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM0__60_carry__0_i_9__2_n_0),
        .I5(PSUM0__60_carry__0_i_10__2_n_0),
        .O(PSUM0__60_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM0__60_carry__0_i_2
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[18]),
        .I2(PSUM0__60_carry__0_i_11_n_0),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM0__60_carry__0_i_2__0
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[2]),
        .I2(PSUM0__60_carry__0_i_11__0_n_0),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM0__60_carry__0_i_2__1
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[18]),
        .I2(PSUM0__60_carry__0_i_11__1_n_0),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM0__60_carry__0_i_2__2
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[2]),
        .I2(PSUM0__60_carry__0_i_11__2_n_0),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM0__60_carry__0_i_3
       (.I0(PSUM0__60_carry__0_i_11_n_0),
        .I1(ALU_DIN2[22]),
        .I2(ALU_DIN1[18]),
        .I3(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ),
        .I5(ALU_DIN1[17]),
        .O(PSUM0__60_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM0__60_carry__0_i_3__0
       (.I0(PSUM0__60_carry__0_i_11__0_n_0),
        .I1(ALU_DIN2[22]),
        .I2(ALU_DIN1[2]),
        .I3(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ),
        .I5(ALU_DIN1[1]),
        .O(PSUM0__60_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM0__60_carry__0_i_3__1
       (.I0(PSUM0__60_carry__0_i_11__1_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[18]),
        .I3(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ),
        .I5(ALU_DIN1[17]),
        .O(PSUM0__60_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM0__60_carry__0_i_3__2
       (.I0(PSUM0__60_carry__0_i_11__2_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[2]),
        .I3(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ),
        .I5(ALU_DIN1[1]),
        .O(PSUM0__60_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM0__60_carry__0_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_7 ),
        .I2(ALU_DIN1[16]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM0__60_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM0__60_carry__0_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_7 ),
        .I2(ALU_DIN1[0]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM0__60_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM0__60_carry__0_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_7 ),
        .I2(ALU_DIN1[16]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM0__60_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM0__60_carry__0_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_7 ),
        .I2(ALU_DIN1[0]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM0__60_carry__0_i_4__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_5
       (.I0(PSUM0__60_carry__0_i_1_n_0),
        .I1(PSUM0__60_carry__0_i_12_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM0__60_carry__0_i_13_n_0),
        .O(PSUM0__60_carry__0_i_5_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_5__0
       (.I0(PSUM0__60_carry__0_i_1__0_n_0),
        .I1(PSUM0__60_carry__0_i_12__0_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM0__60_carry__0_i_13__0_n_0),
        .O(PSUM0__60_carry__0_i_5__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_5__1
       (.I0(PSUM0__60_carry__0_i_1__1_n_0),
        .I1(PSUM0__60_carry__0_i_12__1_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM0__60_carry__0_i_13__1_n_0),
        .O(PSUM0__60_carry__0_i_5__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_5__2
       (.I0(PSUM0__60_carry__0_i_1__2_n_0),
        .I1(PSUM0__60_carry__0_i_12__2_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM0__60_carry__0_i_13__2_n_0),
        .O(PSUM0__60_carry__0_i_5__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_6
       (.I0(PSUM0__60_carry__0_i_2_n_0),
        .I1(PSUM0__60_carry__0_i_9_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM0__60_carry__0_i_10_n_0),
        .O(PSUM0__60_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_6__0
       (.I0(PSUM0__60_carry__0_i_2__0_n_0),
        .I1(PSUM0__60_carry__0_i_9__0_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM0__60_carry__0_i_10__0_n_0),
        .O(PSUM0__60_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_6__1
       (.I0(PSUM0__60_carry__0_i_2__1_n_0),
        .I1(PSUM0__60_carry__0_i_9__1_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM0__60_carry__0_i_10__1_n_0),
        .O(PSUM0__60_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM0__60_carry__0_i_6__2
       (.I0(PSUM0__60_carry__0_i_2__2_n_0),
        .I1(PSUM0__60_carry__0_i_9__2_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM0__60_carry__0_i_10__2_n_0),
        .O(PSUM0__60_carry__0_i_6__2_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM0__60_carry__0_i_7
       (.I0(PSUM0__60_carry__0_i_14_n_0),
        .I1(ALU_DIN1[16]),
        .I2(ALU_DIN2[23]),
        .I3(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_7 ),
        .O(PSUM0__60_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM0__60_carry__0_i_7__0
       (.I0(PSUM0__60_carry__0_i_14__0_n_0),
        .I1(ALU_DIN1[0]),
        .I2(ALU_DIN2[23]),
        .I3(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_7 ),
        .O(PSUM0__60_carry__0_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM0__60_carry__0_i_7__1
       (.I0(PSUM0__60_carry__0_i_14__1_n_0),
        .I1(ALU_DIN1[16]),
        .I2(ALU_DIN2[7]),
        .I3(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_7 ),
        .O(PSUM0__60_carry__0_i_7__1_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM0__60_carry__0_i_7__2
       (.I0(PSUM0__60_carry__0_i_14__2_n_0),
        .I1(ALU_DIN1[0]),
        .I2(ALU_DIN2[7]),
        .I3(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_7 ),
        .O(PSUM0__60_carry__0_i_7__2_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM0__60_carry__0_i_8
       (.I0(PSUM0__60_carry__0_i_15_n_0),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[22]),
        .I3(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_8_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM0__60_carry__0_i_8__0
       (.I0(PSUM0__60_carry__0_i_15__0_n_0),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[22]),
        .I3(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM0__60_carry__0_i_8__1
       (.I0(PSUM0__60_carry__0_i_15__1_n_0),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[6]),
        .I3(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM0__60_carry__0_i_8__2
       (.I0(PSUM0__60_carry__0_i_15__2_n_0),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[6]),
        .I3(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ),
        .O(PSUM0__60_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_9
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[18]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_6 ),
        .O(PSUM0__60_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_9__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[2]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_6 ),
        .O(PSUM0__60_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_9__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[18]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_6 ),
        .O(PSUM0__60_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM0__60_carry__0_i_9__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[2]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_6 ),
        .O(PSUM0__60_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_1
       (.I0(PSUM0__60_carry__1_i_9_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_6 ),
        .I5(ALU_DIN1[21]),
        .O(PSUM0__60_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_10
       (.I0(EX_RF_RD1[6]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[132]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM0__60_carry__1_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_10__0
       (.I0(EX_RF_RD1[22]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[148]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM0__60_carry__1_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM0__60_carry__1_i_10__1
       (.I0(ID_EX_Q[148]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[22]),
        .I3(ID_EX_Q[101]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[22]),
        .O(PSUM0__60_carry__1_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM0__60_carry__1_i_10__2
       (.I0(ID_EX_Q[132]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[6]),
        .I3(ID_EX_Q[85]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[6]),
        .O(PSUM0__60_carry__1_i_10__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__1_i_11
       (.I0(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_1 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[19]),
        .O(PSUM0__60_carry__1_i_11_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__1_i_11__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_1 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[3]),
        .O(PSUM0__60_carry__1_i_11__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__1_i_11__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_1 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[19]),
        .O(PSUM0__60_carry__1_i_11__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM0__60_carry__1_i_11__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_1 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[3]),
        .O(PSUM0__60_carry__1_i_11__2_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_12
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[21]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_12_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_12__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[5]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_12__0_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_12__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[21]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_12__1_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_12__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[5]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_12__2_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM0__60_carry__1_i_13
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[22]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM0__60_carry__1_i_13__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[6]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_13__0_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM0__60_carry__1_i_13__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[22]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_13__1_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM0__60_carry__1_i_13__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[6]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_13__2_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_14
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[20]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_7 ),
        .O(PSUM0__60_carry__1_i_14_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_14__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[4]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_7 ),
        .O(PSUM0__60_carry__1_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_14__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[20]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_7 ),
        .O(PSUM0__60_carry__1_i_14__1_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM0__60_carry__1_i_14__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[4]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_7 ),
        .O(PSUM0__60_carry__1_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_15
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM0__60_carry__1_i_15_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_15__0
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM0__60_carry__1_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_15__1
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM0__60_carry__1_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_15__2
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM0__60_carry__1_i_15__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_1__0
       (.I0(PSUM0__60_carry__1_i_9__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_6 ),
        .I5(ALU_DIN1[5]),
        .O(PSUM0__60_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_1__1
       (.I0(PSUM0__60_carry__1_i_9__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_6 ),
        .I5(ALU_DIN1[21]),
        .O(PSUM0__60_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_1__2
       (.I0(PSUM0__60_carry__1_i_9__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_6 ),
        .I5(ALU_DIN1[5]),
        .O(PSUM0__60_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_2
       (.I0(PSUM0__60_carry__1_i_10__1_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_7 ),
        .I5(ALU_DIN1[20]),
        .O(PSUM0__60_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_2__0
       (.I0(PSUM0__60_carry__1_i_10__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_7 ),
        .I5(ALU_DIN1[4]),
        .O(PSUM0__60_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_2__1
       (.I0(PSUM0__60_carry__1_i_10_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_7 ),
        .I5(ALU_DIN1[4]),
        .O(PSUM0__60_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM0__60_carry__1_i_2__2
       (.I0(PSUM0__60_carry__1_i_10__0_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_7 ),
        .I5(ALU_DIN1[20]),
        .O(PSUM0__60_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM0__60_carry__1_i_3
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[21]),
        .I2(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_7 ),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[23]),
        .I5(PSUM0__60_carry__1_i_11_n_0),
        .O(PSUM0__60_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM0__60_carry__1_i_3__0
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[5]),
        .I2(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_7 ),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[23]),
        .I5(PSUM0__60_carry__1_i_11__0_n_0),
        .O(PSUM0__60_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM0__60_carry__1_i_3__1
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[21]),
        .I2(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_7 ),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[7]),
        .I5(PSUM0__60_carry__1_i_11__1_n_0),
        .O(PSUM0__60_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM0__60_carry__1_i_3__2
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[5]),
        .I2(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_7 ),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[7]),
        .I5(PSUM0__60_carry__1_i_11__2_n_0),
        .O(PSUM0__60_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__1_i_4
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM0__60_carry__0_i_12_n_0),
        .I5(PSUM0__60_carry__0_i_13_n_0),
        .O(PSUM0__60_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__1_i_4__0
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM0__60_carry__0_i_12__0_n_0),
        .I5(PSUM0__60_carry__0_i_13__0_n_0),
        .O(PSUM0__60_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__1_i_4__1
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM0__60_carry__0_i_12__1_n_0),
        .I5(PSUM0__60_carry__0_i_13__1_n_0),
        .O(PSUM0__60_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM0__60_carry__1_i_4__2
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM0__60_carry__0_i_12__2_n_0),
        .I5(PSUM0__60_carry__0_i_13__2_n_0),
        .O(PSUM0__60_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM0__60_carry__1_i_5
       (.I0(PSUM0__60_carry__1_i_12_n_0),
        .I1(ALU_DIN2[22]),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[22]),
        .I5(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_5_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM0__60_carry__1_i_5__0
       (.I0(PSUM0__60_carry__1_i_12__2_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[7]),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[6]),
        .I5(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM0__60_carry__1_i_5__1
       (.I0(PSUM0__60_carry__1_i_12__0_n_0),
        .I1(ALU_DIN2[22]),
        .I2(ALU_DIN1[7]),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[6]),
        .I5(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM0__60_carry__1_i_5__2
       (.I0(PSUM0__60_carry__1_i_12__1_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[22]),
        .I5(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_1 ),
        .O(PSUM0__60_carry__1_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM0__60_carry__1_i_6
       (.I0(PSUM0__60_carry__1_i_2_n_0),
        .I1(PSUM0__60_carry__1_i_13_n_0),
        .I2(PSUM0__60_carry__1_i_9_n_0),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[21]),
        .I5(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_6_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM0__60_carry__1_i_6__0
       (.I0(PSUM0__60_carry__1_i_2__0_n_0),
        .I1(PSUM0__60_carry__1_i_13__2_n_0),
        .I2(PSUM0__60_carry__1_i_9__2_n_0),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[5]),
        .I5(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM0__60_carry__1_i_6__1
       (.I0(PSUM0__60_carry__1_i_2__1_n_0),
        .I1(PSUM0__60_carry__1_i_13__0_n_0),
        .I2(PSUM0__60_carry__1_i_9__0_n_0),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[5]),
        .I5(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM0__60_carry__1_i_6__2
       (.I0(PSUM0__60_carry__1_i_2__2_n_0),
        .I1(PSUM0__60_carry__1_i_13__1_n_0),
        .I2(PSUM0__60_carry__1_i_9__1_n_0),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[21]),
        .I5(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_6 ),
        .O(PSUM0__60_carry__1_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM0__60_carry__1_i_7
       (.I0(PSUM0__60_carry__1_i_3_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[23]),
        .I4(PSUM0__60_carry__1_i_10__1_n_0),
        .I5(PSUM0__60_carry__1_i_14_n_0),
        .O(PSUM0__60_carry__1_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM0__60_carry__1_i_7__0
       (.I0(PSUM0__60_carry__1_i_3__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[7]),
        .I4(PSUM0__60_carry__1_i_10__2_n_0),
        .I5(PSUM0__60_carry__1_i_14__2_n_0),
        .O(PSUM0__60_carry__1_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM0__60_carry__1_i_7__1
       (.I0(PSUM0__60_carry__1_i_3__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[23]),
        .I4(PSUM0__60_carry__1_i_10_n_0),
        .I5(PSUM0__60_carry__1_i_14__0_n_0),
        .O(PSUM0__60_carry__1_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM0__60_carry__1_i_7__2
       (.I0(PSUM0__60_carry__1_i_3__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[7]),
        .I4(PSUM0__60_carry__1_i_10__0_n_0),
        .I5(PSUM0__60_carry__1_i_14__1_n_0),
        .O(PSUM0__60_carry__1_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM0__60_carry__1_i_8
       (.I0(PSUM0__60_carry__1_i_4_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_7 ),
        .I2(ALU_DIN1[20]),
        .I3(ALU_DIN2[23]),
        .I4(PSUM0__60_carry__1_i_15_n_0),
        .I5(PSUM0__60_carry__1_i_11_n_0),
        .O(PSUM0__60_carry__1_i_8_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM0__60_carry__1_i_8__0
       (.I0(PSUM0__60_carry__1_i_4__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_7 ),
        .I2(ALU_DIN1[4]),
        .I3(ALU_DIN2[23]),
        .I4(PSUM0__60_carry__1_i_15__0_n_0),
        .I5(PSUM0__60_carry__1_i_11__0_n_0),
        .O(PSUM0__60_carry__1_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM0__60_carry__1_i_8__1
       (.I0(PSUM0__60_carry__1_i_4__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_7 ),
        .I2(ALU_DIN1[20]),
        .I3(ALU_DIN2[7]),
        .I4(PSUM0__60_carry__1_i_15__1_n_0),
        .I5(PSUM0__60_carry__1_i_11__1_n_0),
        .O(PSUM0__60_carry__1_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM0__60_carry__1_i_8__2
       (.I0(PSUM0__60_carry__1_i_4__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_7 ),
        .I2(ALU_DIN1[4]),
        .I3(ALU_DIN2[7]),
        .I4(PSUM0__60_carry__1_i_15__2_n_0),
        .I5(PSUM0__60_carry__1_i_11__2_n_0),
        .O(PSUM0__60_carry__1_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_9
       (.I0(EX_RF_RD1[23]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[149]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM0__60_carry__1_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_9__0
       (.I0(EX_RF_RD1[7]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[133]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM0__60_carry__1_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_9__1
       (.I0(EX_RF_RD1[23]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[149]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM0__60_carry__1_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM0__60_carry__1_i_9__2
       (.I0(EX_RF_RD1[7]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[133]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM0__60_carry__1_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM0__60_carry__2_i_1
       (.I0(ALU_DIN1[23]),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM0__60_carry__2_i_1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM0__60_carry__2_i_1__0
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM0__60_carry__2_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM0__60_carry__2_i_1__1
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM0__60_carry__2_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM0__60_carry__2_i_1__2
       (.I0(ALU_DIN1[23]),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM0__60_carry__2_i_1__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_1
       (.I0(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ),
        .O(PSUM0__60_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_1__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ),
        .O(PSUM0__60_carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_1__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ),
        .O(PSUM0__60_carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_1__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ),
        .O(PSUM0__60_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM0__60_carry_i_2
       (.I0(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ),
        .I2(ID_EX_Q[101]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[22]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__60_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM0__60_carry_i_2__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ),
        .I2(ID_EX_Q[101]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[22]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__60_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM0__60_carry_i_2__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ),
        .I2(ID_EX_Q[85]),
        .I3(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I4(EX_RF_RD2[6]),
        .I5(ALU_DIN1[16]),
        .O(PSUM0__60_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM0__60_carry_i_2__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ),
        .I2(ID_EX_Q[85]),
        .I3(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I4(EX_RF_RD2[6]),
        .I5(ALU_DIN1[0]),
        .O(PSUM0__60_carry_i_2__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_3
       (.I0(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_5 ),
        .O(PSUM0__60_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_3__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_5 ),
        .O(PSUM0__60_carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_3__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_5 ),
        .O(PSUM0__60_carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_3__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_5 ),
        .O(PSUM0__60_carry_i_3__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_6 ),
        .O(PSUM0__60_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_6 ),
        .O(PSUM0__60_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_6 ),
        .O(PSUM0__60_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_6 ),
        .O(PSUM0__60_carry_i_4__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_5
       (.I0(\custom_alu/mult/mult16_3/PSUM0__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_7 ),
        .O(PSUM0__60_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_5__0
       (.I0(\custom_alu/mult/mult16_2/PSUM0__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_7 ),
        .O(PSUM0__60_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_5__1
       (.I0(\custom_alu/mult/mult16_1/PSUM0__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_7 ),
        .O(PSUM0__60_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM0__60_carry_i_5__2
       (.I0(\custom_alu/mult/mult16_0/PSUM0__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_7 ),
        .O(PSUM0__60_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_1
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[30]),
        .O(PSUM1__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_10
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM1__0_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_10__0
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM1__0_carry__0_i_10__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_10__1
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(ALU_DIN2[2]),
        .O(PSUM1__0_carry__0_i_10__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1__0_carry__0_i_10__2
       (.I0(ID_EX_Q[157]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[31]),
        .O(ALU_DIN1[31]));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_11
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM1__0_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_11__0
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[17]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[96]),
        .O(PSUM1__0_carry__0_i_11__0_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_11__1
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(ALU_DIN2[2]),
        .O(PSUM1__0_carry__0_i_11__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_11__2
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(ALU_DIN2[1]),
        .O(PSUM1__0_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_12
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM1__0_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_12__0
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[136]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM1__0_carry__0_i_12__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_12__1
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(ALU_DIN2[2]),
        .O(PSUM1__0_carry__0_i_12__1_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_12__2
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[136]),
        .I3(ALU_DIN2[2]),
        .O(PSUM1__0_carry__0_i_12__2_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_13
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(ALU_DIN2[2]),
        .O(PSUM1__0_carry__0_i_13_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_1__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[14]),
        .O(PSUM1__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_1__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[30]),
        .O(PSUM1__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_1__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[14]),
        .O(PSUM1__0_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_2
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[29]),
        .O(PSUM1__0_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_2__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[13]),
        .O(PSUM1__0_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_2__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[29]),
        .O(PSUM1__0_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_2__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[13]),
        .O(PSUM1__0_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_3
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[28]),
        .O(PSUM1__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_3__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[12]),
        .O(PSUM1__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_3__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[28]),
        .O(PSUM1__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_3__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[12]),
        .O(PSUM1__0_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_4
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[27]),
        .O(PSUM1__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_4__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[11]),
        .O(PSUM1__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_4__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[27]),
        .O(PSUM1__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__0_i_4__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[11]),
        .O(PSUM1__0_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_5
       (.I0(PSUM1__0_carry__0_i_1_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM1__0_carry__0_i_9_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_5__0
       (.I0(PSUM1__0_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM1__0_carry__0_i_9__0_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_5__1
       (.I0(PSUM1__0_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM1__0_carry__0_i_9__1_n_0),
        .I4(ALU_DIN1[31]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_5__2
       (.I0(PSUM1__0_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM1__0_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_6
       (.I0(PSUM1__0_carry__0_i_2_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM1__0_carry__0_i_10_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_6__0
       (.I0(PSUM1__0_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM1__0_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_6__1
       (.I0(PSUM1__0_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM1__0_carry__0_i_11__1_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_6__2
       (.I0(PSUM1__0_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM1__0_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_7
       (.I0(PSUM1__0_carry__0_i_3_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM1__0_carry__0_i_11_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM1__0_carry__0_i_7__0
       (.I0(PSUM1__0_carry__0_i_3__0_n_0),
        .I1(PSUM1__0_carry__0_i_11__0_n_0),
        .I2(ALU_DIN2[18]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_7__1
       (.I0(PSUM1__0_carry__0_i_3__1_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM1__0_carry__0_i_12__1_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM1__0_carry__0_i_7__2
       (.I0(PSUM1__0_carry__0_i_3__2_n_0),
        .I1(PSUM1__0_carry__0_i_11__2_n_0),
        .I2(ALU_DIN2[2]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_8
       (.I0(PSUM1__0_carry__0_i_4_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM1__0_carry__0_i_12_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_8__0
       (.I0(PSUM1__0_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[17]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM1__0_carry__0_i_12__0_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_8__1
       (.I0(PSUM1__0_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM1__0_carry__0_i_13_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__0_carry__0_i_8__2
       (.I0(PSUM1__0_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[1]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM1__0_carry__0_i_12__2_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_9
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM1__0_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry__0_i_9__0
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[18]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[97]),
        .O(PSUM1__0_carry__0_i_9__0_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_9__1
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(ALU_DIN2[2]),
        .O(PSUM1__0_carry__0_i_9__1_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry__0_i_9__2
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(ALU_DIN2[2]),
        .O(PSUM1__0_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM1__0_carry__1_i_1
       (.I0(ID_EX_Q[97]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[18]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[17]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM1__0_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM1__0_carry__1_i_1__0
       (.I0(ID_EX_Q[97]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[18]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[17]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__0_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM1__0_carry__1_i_1__1
       (.I0(ALU_DIN2[2]),
        .I1(ID_EX_Q[156]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[30]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[31]),
        .O(PSUM1__0_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM1__0_carry__1_i_1__2
       (.I0(ALU_DIN2[2]),
        .I1(ID_EX_Q[140]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[14]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__0_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__1_i_2
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[16]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM1__0_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__1_i_2__0
       (.I0(ALU_DIN2[18]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[17]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__0_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__1_i_2__1
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[31]),
        .O(PSUM1__0_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__0_carry__1_i_2__2
       (.I0(ALU_DIN2[2]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[1]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__0_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM1__0_carry__1_i_3
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[96]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[18]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM1__0_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM1__0_carry__1_i_3__0
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[96]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[18]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__0_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM1__0_carry__1_i_3__1
       (.I0(ALU_DIN2[1]),
        .I1(EX_RF_RD1[30]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[156]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[31]),
        .O(PSUM1__0_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM1__0_carry__1_i_3__2
       (.I0(ALU_DIN2[1]),
        .I1(EX_RF_RD1[14]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[140]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__0_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__0_carry__1_i_4
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[18]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[17]),
        .O(PSUM1__0_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__0_carry__1_i_4__0
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[18]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[17]),
        .O(PSUM1__0_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__0_carry__1_i_4__1
       (.I0(ALU_DIN2[0]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[2]),
        .I4(ALU_DIN1[31]),
        .I5(ALU_DIN2[1]),
        .O(PSUM1__0_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__0_carry__1_i_4__2
       (.I0(ALU_DIN2[0]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[2]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[1]),
        .O(PSUM1__0_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_1
       (.I0(ALU_DIN2[17]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[18]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_1__0
       (.I0(ALU_DIN2[17]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[18]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[16]),
        .O(PSUM1__0_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_1__1
       (.I0(ALU_DIN2[1]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[2]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_1__2
       (.I0(ALU_DIN2[1]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[2]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[0]),
        .O(PSUM1__0_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM1__0_carry_i_2
       (.I0(ID_EX_Q[96]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[17]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[18]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__0_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM1__0_carry_i_2__0
       (.I0(ID_EX_Q[96]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[17]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[18]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__0_carry_i_2__1
       (.I0(ALU_DIN2[1]),
        .I1(ID_EX_Q[151]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[25]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__0_carry_i_2__2
       (.I0(ALU_DIN2[1]),
        .I1(ID_EX_Q[135]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[9]),
        .I4(ALU_DIN2[2]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__0_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM1__0_carry_i_3
       (.I0(ID_EX_Q[95]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[16]),
        .I3(ID_EX_Q[151]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[25]),
        .O(PSUM1__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM1__0_carry_i_3__0
       (.I0(ID_EX_Q[95]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[16]),
        .I3(ID_EX_Q[135]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[9]),
        .O(PSUM1__0_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM1__0_carry_i_3__1
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[151]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[25]),
        .O(PSUM1__0_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM1__0_carry_i_3__2
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[135]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[9]),
        .O(PSUM1__0_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__0_carry_i_4
       (.I0(ALU_DIN1[26]),
        .I1(PSUM1__0_carry_i_8_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[18]),
        .O(PSUM1__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__0_carry_i_4__0
       (.I0(ALU_DIN1[10]),
        .I1(PSUM1__0_carry_i_8__0_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[18]),
        .O(PSUM1__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__0_carry_i_4__1
       (.I0(ALU_DIN1[26]),
        .I1(PSUM1__0_carry_i_8__1_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[2]),
        .O(PSUM1__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__0_carry_i_4__2
       (.I0(ALU_DIN1[10]),
        .I1(PSUM1__0_carry_i_8__2_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[2]),
        .O(PSUM1__0_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_5
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[18]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[26]),
        .O(PSUM1__0_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_5__0
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[18]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[17]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[10]),
        .O(PSUM1__0_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_5__1
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[26]),
        .O(PSUM1__0_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__0_carry_i_5__2
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[2]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[10]),
        .O(PSUM1__0_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM1__0_carry_i_6
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[25]),
        .I2(ID_EX_Q[96]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[17]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__0_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM1__0_carry_i_6__0
       (.I0(ALU_DIN2[16]),
        .I1(ALU_DIN1[9]),
        .I2(ID_EX_Q[96]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[17]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__0_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__0_carry_i_6__1
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[151]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[25]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__0_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__0_carry_i_6__2
       (.I0(ALU_DIN2[0]),
        .I1(ID_EX_Q[135]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[9]),
        .I4(ALU_DIN2[1]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__0_carry_i_6__2_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    PSUM1__0_carry_i_7
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(ALU_DIN2[0]),
        .O(PSUM1__0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM1__0_carry_i_7__0
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM1__0_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    PSUM1__0_carry_i_7__1
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(ALU_DIN2[0]),
        .O(PSUM1__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM1__0_carry_i_7__2
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM1__0_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry_i_8
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM1__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__0_carry_i_8__0
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(EX_RF_RD2[16]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[95]),
        .O(PSUM1__0_carry_i_8__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry_i_8__1
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(ALU_DIN2[0]),
        .O(PSUM1__0_carry_i_8__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__0_carry_i_8__2
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(ALU_DIN2[0]),
        .O(PSUM1__0_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_1
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[30]),
        .O(PSUM1__30_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_10
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM1__30_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_10__0
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM1__30_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_10__1
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_10__2
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_11
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM1__30_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_11__0
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[20]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[99]),
        .O(PSUM1__30_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_11__1
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_11__2
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_12
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM1__30_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_12__0
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[136]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM1__30_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_12__1
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_12__2
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[136]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_1__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[14]),
        .O(PSUM1__30_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_1__1
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[30]),
        .O(PSUM1__30_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_1__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[14]),
        .O(PSUM1__30_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_2
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[29]),
        .O(PSUM1__30_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_2__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[13]),
        .O(PSUM1__30_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_2__1
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[29]),
        .O(PSUM1__30_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_2__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[13]),
        .O(PSUM1__30_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_3
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[28]),
        .O(PSUM1__30_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_3__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[12]),
        .O(PSUM1__30_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_3__1
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[28]),
        .O(PSUM1__30_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_3__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[12]),
        .O(PSUM1__30_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_4
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[27]),
        .O(PSUM1__30_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_4__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[11]),
        .O(PSUM1__30_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_4__1
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[27]),
        .O(PSUM1__30_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__0_i_4__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[11]),
        .O(PSUM1__30_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_5
       (.I0(PSUM1__30_carry__0_i_1_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM1__30_carry__0_i_9_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_5__0
       (.I0(PSUM1__30_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM1__30_carry__0_i_9__0_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_5__1
       (.I0(PSUM1__30_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM1__30_carry__0_i_9__1_n_0),
        .I4(ALU_DIN1[31]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_5__2
       (.I0(PSUM1__30_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM1__30_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_6
       (.I0(PSUM1__30_carry__0_i_2_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM1__30_carry__0_i_10_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_6__0
       (.I0(PSUM1__30_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM1__30_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_6__1
       (.I0(PSUM1__30_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM1__30_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_6__2
       (.I0(PSUM1__30_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM1__30_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_7
       (.I0(PSUM1__30_carry__0_i_3_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM1__30_carry__0_i_11_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM1__30_carry__0_i_7__0
       (.I0(PSUM1__30_carry__0_i_3__0_n_0),
        .I1(PSUM1__30_carry__0_i_11__0_n_0),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_7__1
       (.I0(PSUM1__30_carry__0_i_3__1_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM1__30_carry__0_i_11__1_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_7__2
       (.I0(PSUM1__30_carry__0_i_3__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[12]),
        .I3(PSUM1__30_carry__0_i_11__2_n_0),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_8
       (.I0(PSUM1__30_carry__0_i_4_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM1__30_carry__0_i_12_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_8__0
       (.I0(PSUM1__30_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[20]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM1__30_carry__0_i_12__0_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_8__1
       (.I0(PSUM1__30_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM1__30_carry__0_i_12__1_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM1__30_carry__0_i_8__2
       (.I0(PSUM1__30_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[4]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM1__30_carry__0_i_12__2_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_9
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM1__30_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_9__0
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[21]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[100]),
        .O(PSUM1__30_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_9__1
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry__0_i_9__2
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[5]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[84]),
        .O(PSUM1__30_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM1__30_carry__1_i_1
       (.I0(ID_EX_Q[100]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[21]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[20]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM1__30_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM1__30_carry__1_i_1__0
       (.I0(ID_EX_Q[100]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[21]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[20]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__30_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM1__30_carry__1_i_1__1
       (.I0(ALU_DIN2[5]),
        .I1(ID_EX_Q[156]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[30]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[31]),
        .O(PSUM1__30_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8A80000000000000)) 
    PSUM1__30_carry__1_i_1__2
       (.I0(ALU_DIN2[5]),
        .I1(ID_EX_Q[140]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[14]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__30_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__1_i_2
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[19]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM1__30_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__1_i_2__0
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[20]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__30_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__1_i_2__1
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[31]),
        .O(PSUM1__30_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM1__30_carry__1_i_2__2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[4]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__30_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM1__30_carry__1_i_3
       (.I0(EX_RF_RD2[20]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[99]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[21]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM1__30_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM1__30_carry__1_i_3__0
       (.I0(EX_RF_RD2[20]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[99]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[21]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__30_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM1__30_carry__1_i_3__1
       (.I0(ALU_DIN2[4]),
        .I1(EX_RF_RD1[30]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[156]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[31]),
        .O(PSUM1__30_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h57F7000000000000)) 
    PSUM1__30_carry__1_i_3__2
       (.I0(ALU_DIN2[4]),
        .I1(EX_RF_RD1[14]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[140]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[15]),
        .O(PSUM1__30_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__30_carry__1_i_4
       (.I0(ALU_DIN2[19]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[21]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[20]),
        .O(PSUM1__30_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__30_carry__1_i_4__0
       (.I0(ALU_DIN2[19]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[21]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[20]),
        .O(PSUM1__30_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__30_carry__1_i_4__1
       (.I0(ALU_DIN2[3]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[31]),
        .I5(ALU_DIN2[4]),
        .O(PSUM1__30_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM1__30_carry__1_i_4__2
       (.I0(ALU_DIN2[3]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[5]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[4]),
        .O(PSUM1__30_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_1
       (.I0(ALU_DIN2[20]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_1__0
       (.I0(ALU_DIN2[20]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[21]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[19]),
        .O(PSUM1__30_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_1__1
       (.I0(ALU_DIN2[4]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_1__2
       (.I0(ALU_DIN2[4]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[5]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[3]),
        .O(PSUM1__30_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM1__30_carry_i_2
       (.I0(ID_EX_Q[99]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[20]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[21]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__30_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM1__30_carry_i_2__0
       (.I0(ID_EX_Q[99]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[20]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[21]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__30_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__30_carry_i_2__1
       (.I0(ALU_DIN2[4]),
        .I1(ID_EX_Q[151]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[25]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__30_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__30_carry_i_2__2
       (.I0(ALU_DIN2[4]),
        .I1(ID_EX_Q[135]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[9]),
        .I4(ALU_DIN2[5]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__30_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM1__30_carry_i_3
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ID_EX_Q[151]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[25]),
        .O(PSUM1__30_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM1__30_carry_i_3__0
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ID_EX_Q[135]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[9]),
        .O(PSUM1__30_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM1__30_carry_i_3__1
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[151]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[25]),
        .O(PSUM1__30_carry_i_3__1_n_0));
  LUT4 #(
    .INIT(16'h8A80)) 
    PSUM1__30_carry_i_3__2
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[135]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[9]),
        .O(PSUM1__30_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__30_carry_i_4
       (.I0(ALU_DIN1[26]),
        .I1(PSUM1__30_carry_i_8_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[21]),
        .O(PSUM1__30_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__30_carry_i_4__0
       (.I0(ALU_DIN1[10]),
        .I1(PSUM1__30_carry_i_8__0_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[21]),
        .O(PSUM1__30_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__30_carry_i_4__1
       (.I0(ALU_DIN1[26]),
        .I1(PSUM1__30_carry_i_8__1_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[5]),
        .O(PSUM1__30_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM1__30_carry_i_4__2
       (.I0(ALU_DIN1[10]),
        .I1(PSUM1__30_carry_i_8__2_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[5]),
        .O(PSUM1__30_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_5
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[21]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[26]),
        .O(PSUM1__30_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_5__0
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[21]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[20]),
        .I4(ALU_DIN2[19]),
        .I5(ALU_DIN1[10]),
        .O(PSUM1__30_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_5__1
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[5]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[26]),
        .O(PSUM1__30_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM1__30_carry_i_5__2
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[5]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[4]),
        .I4(ALU_DIN2[3]),
        .I5(ALU_DIN1[10]),
        .O(PSUM1__30_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM1__30_carry_i_6
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[20]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__30_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM1__30_carry_i_6__0
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[20]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__30_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__30_carry_i_6__1
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[151]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[25]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__30_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h757F8A808A808A80)) 
    PSUM1__30_carry_i_6__2
       (.I0(ALU_DIN2[3]),
        .I1(ID_EX_Q[135]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[9]),
        .I4(ALU_DIN2[4]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__30_carry_i_6__2_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    PSUM1__30_carry_i_7
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(ALU_DIN2[3]),
        .O(PSUM1__30_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM1__30_carry_i_7__0
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM1__30_carry_i_7__0_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    PSUM1__30_carry_i_7__1
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(ALU_DIN2[3]),
        .O(PSUM1__30_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM1__30_carry_i_7__2
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM1__30_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry_i_8
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM1__30_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__30_carry_i_8__0
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(EX_RF_RD2[19]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[98]),
        .O(PSUM1__30_carry_i_8__0_n_0));
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__30_carry_i_8__1
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(ALU_DIN2[3]),
        .O(PSUM1__30_carry_i_8__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    PSUM1__30_carry_i_8__2
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(ALU_DIN2[3]),
        .O(PSUM1__30_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__0_i_1
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM1__60_carry__0_i_9_n_0),
        .I5(PSUM1__60_carry__0_i_10_n_0),
        .O(PSUM1__60_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_10
       (.I0(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_7 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[25]),
        .O(PSUM1__60_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_10__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_7 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[9]),
        .O(PSUM1__60_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_10__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_7 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[25]),
        .O(PSUM1__60_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_10__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_7 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[9]),
        .O(PSUM1__60_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_11
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_7 ),
        .O(PSUM1__60_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_11__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_7 ),
        .O(PSUM1__60_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_11__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_7 ),
        .O(PSUM1__60_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_11__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_7 ),
        .O(PSUM1__60_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_12
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[27]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_1 ),
        .O(PSUM1__60_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_12__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[11]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_1 ),
        .O(PSUM1__60_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_12__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[27]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_1 ),
        .O(PSUM1__60_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_12__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[11]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_1 ),
        .O(PSUM1__60_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_13
       (.I0(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_6 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[26]),
        .O(PSUM1__60_carry__0_i_13_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_13__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_6 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[10]),
        .O(PSUM1__60_carry__0_i_13__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_13__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_6 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[26]),
        .O(PSUM1__60_carry__0_i_13__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__0_i_13__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_6 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[10]),
        .O(PSUM1__60_carry__0_i_13__2_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM1__60_carry__0_i_14
       (.I0(ALU_DIN1[25]),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[22]),
        .I5(PSUM1__60_carry__0_i_11_n_0),
        .O(PSUM1__60_carry__0_i_14_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM1__60_carry__0_i_14__0
       (.I0(ALU_DIN1[9]),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[22]),
        .I5(PSUM1__60_carry__0_i_11__0_n_0),
        .O(PSUM1__60_carry__0_i_14__0_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM1__60_carry__0_i_14__1
       (.I0(ALU_DIN1[25]),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[6]),
        .I5(PSUM1__60_carry__0_i_11__1_n_0),
        .O(PSUM1__60_carry__0_i_14__1_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM1__60_carry__0_i_14__2
       (.I0(ALU_DIN1[9]),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[6]),
        .I5(PSUM1__60_carry__0_i_11__2_n_0),
        .O(PSUM1__60_carry__0_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_15
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[24]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_4 ),
        .O(PSUM1__60_carry__0_i_15_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_15__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[8]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_4 ),
        .O(PSUM1__60_carry__0_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_15__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[24]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_4 ),
        .O(PSUM1__60_carry__0_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_15__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[8]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_4 ),
        .O(PSUM1__60_carry__0_i_15__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__0_i_1__0
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM1__60_carry__0_i_9__0_n_0),
        .I5(PSUM1__60_carry__0_i_10__0_n_0),
        .O(PSUM1__60_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__0_i_1__1
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM1__60_carry__0_i_9__1_n_0),
        .I5(PSUM1__60_carry__0_i_10__1_n_0),
        .O(PSUM1__60_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__0_i_1__2
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM1__60_carry__0_i_9__2_n_0),
        .I5(PSUM1__60_carry__0_i_10__2_n_0),
        .O(PSUM1__60_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM1__60_carry__0_i_2
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[26]),
        .I2(PSUM1__60_carry__0_i_11_n_0),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM1__60_carry__0_i_2__0
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[10]),
        .I2(PSUM1__60_carry__0_i_11__0_n_0),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM1__60_carry__0_i_2__1
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[26]),
        .I2(PSUM1__60_carry__0_i_11__1_n_0),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM1__60_carry__0_i_2__2
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[10]),
        .I2(PSUM1__60_carry__0_i_11__2_n_0),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM1__60_carry__0_i_3
       (.I0(PSUM1__60_carry__0_i_11_n_0),
        .I1(ALU_DIN2[22]),
        .I2(ALU_DIN1[26]),
        .I3(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ),
        .I5(ALU_DIN1[25]),
        .O(PSUM1__60_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM1__60_carry__0_i_3__0
       (.I0(PSUM1__60_carry__0_i_11__0_n_0),
        .I1(ALU_DIN2[22]),
        .I2(ALU_DIN1[10]),
        .I3(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ),
        .I5(ALU_DIN1[9]),
        .O(PSUM1__60_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM1__60_carry__0_i_3__1
       (.I0(PSUM1__60_carry__0_i_11__1_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[26]),
        .I3(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ),
        .I5(ALU_DIN1[25]),
        .O(PSUM1__60_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM1__60_carry__0_i_3__2
       (.I0(PSUM1__60_carry__0_i_11__2_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[10]),
        .I3(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ),
        .I5(ALU_DIN1[9]),
        .O(PSUM1__60_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM1__60_carry__0_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_7 ),
        .I2(ALU_DIN1[24]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM1__60_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM1__60_carry__0_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_7 ),
        .I2(ALU_DIN1[8]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM1__60_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM1__60_carry__0_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_7 ),
        .I2(ALU_DIN1[24]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM1__60_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM1__60_carry__0_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_7 ),
        .I2(ALU_DIN1[8]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM1__60_carry__0_i_4__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_5
       (.I0(PSUM1__60_carry__0_i_1_n_0),
        .I1(PSUM1__60_carry__0_i_12_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM1__60_carry__0_i_13_n_0),
        .O(PSUM1__60_carry__0_i_5_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_5__0
       (.I0(PSUM1__60_carry__0_i_1__0_n_0),
        .I1(PSUM1__60_carry__0_i_12__0_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM1__60_carry__0_i_13__0_n_0),
        .O(PSUM1__60_carry__0_i_5__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_5__1
       (.I0(PSUM1__60_carry__0_i_1__1_n_0),
        .I1(PSUM1__60_carry__0_i_12__1_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM1__60_carry__0_i_13__1_n_0),
        .O(PSUM1__60_carry__0_i_5__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_5__2
       (.I0(PSUM1__60_carry__0_i_1__2_n_0),
        .I1(PSUM1__60_carry__0_i_12__2_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM1__60_carry__0_i_13__2_n_0),
        .O(PSUM1__60_carry__0_i_5__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_6
       (.I0(PSUM1__60_carry__0_i_2_n_0),
        .I1(PSUM1__60_carry__0_i_9_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM1__60_carry__0_i_10_n_0),
        .O(PSUM1__60_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_6__0
       (.I0(PSUM1__60_carry__0_i_2__0_n_0),
        .I1(PSUM1__60_carry__0_i_9__0_n_0),
        .I2(ALU_DIN2[22]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM1__60_carry__0_i_10__0_n_0),
        .O(PSUM1__60_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_6__1
       (.I0(PSUM1__60_carry__0_i_2__1_n_0),
        .I1(PSUM1__60_carry__0_i_9__1_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM1__60_carry__0_i_10__1_n_0),
        .O(PSUM1__60_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM1__60_carry__0_i_6__2
       (.I0(PSUM1__60_carry__0_i_2__2_n_0),
        .I1(PSUM1__60_carry__0_i_9__2_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM1__60_carry__0_i_10__2_n_0),
        .O(PSUM1__60_carry__0_i_6__2_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM1__60_carry__0_i_7
       (.I0(PSUM1__60_carry__0_i_14_n_0),
        .I1(ALU_DIN1[24]),
        .I2(ALU_DIN2[23]),
        .I3(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_7 ),
        .O(PSUM1__60_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM1__60_carry__0_i_7__0
       (.I0(PSUM1__60_carry__0_i_14__0_n_0),
        .I1(ALU_DIN1[8]),
        .I2(ALU_DIN2[23]),
        .I3(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_7 ),
        .O(PSUM1__60_carry__0_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM1__60_carry__0_i_7__1
       (.I0(PSUM1__60_carry__0_i_14__1_n_0),
        .I1(ALU_DIN1[24]),
        .I2(ALU_DIN2[7]),
        .I3(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_7 ),
        .O(PSUM1__60_carry__0_i_7__1_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM1__60_carry__0_i_7__2
       (.I0(PSUM1__60_carry__0_i_14__2_n_0),
        .I1(ALU_DIN1[8]),
        .I2(ALU_DIN2[7]),
        .I3(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_7 ),
        .O(PSUM1__60_carry__0_i_7__2_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM1__60_carry__0_i_8
       (.I0(PSUM1__60_carry__0_i_15_n_0),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[22]),
        .I3(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_8_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM1__60_carry__0_i_8__0
       (.I0(PSUM1__60_carry__0_i_15__0_n_0),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[22]),
        .I3(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM1__60_carry__0_i_8__1
       (.I0(PSUM1__60_carry__0_i_15__1_n_0),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[6]),
        .I3(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM1__60_carry__0_i_8__2
       (.I0(PSUM1__60_carry__0_i_15__2_n_0),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[6]),
        .I3(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ),
        .O(PSUM1__60_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_9
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[26]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_6 ),
        .O(PSUM1__60_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_9__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[10]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_6 ),
        .O(PSUM1__60_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_9__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[26]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_6 ),
        .O(PSUM1__60_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM1__60_carry__0_i_9__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[10]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_6 ),
        .O(PSUM1__60_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_1
       (.I0(PSUM1__60_carry__1_i_9_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_6 ),
        .I5(ALU_DIN1[29]),
        .O(PSUM1__60_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_10
       (.I0(EX_RF_RD1[30]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[156]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM1__60_carry__1_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_10__0
       (.I0(EX_RF_RD1[14]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[140]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM1__60_carry__1_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_10__1
       (.I0(EX_RF_RD1[30]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[156]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM1__60_carry__1_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_10__2
       (.I0(EX_RF_RD1[14]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[140]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM1__60_carry__1_i_10__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__1_i_11
       (.I0(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_1 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[27]),
        .O(PSUM1__60_carry__1_i_11_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__1_i_11__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_1 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[23]),
        .I5(ALU_DIN1[11]),
        .O(PSUM1__60_carry__1_i_11__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__1_i_11__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_1 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[27]),
        .O(PSUM1__60_carry__1_i_11__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM1__60_carry__1_i_11__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_1 ),
        .I2(ID_EX_Q[86]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[7]),
        .I5(ALU_DIN1[11]),
        .O(PSUM1__60_carry__1_i_11__2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM1__60_carry__1_i_12
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM1__60_carry__1_i_12__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_12__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM1__60_carry__1_i_12__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_12__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM1__60_carry__1_i_12__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_12__2_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_13
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[30]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_13__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[14]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_13__0_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_13__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[30]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_13__1_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_13__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[14]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_13__2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_14
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_14_n_0));
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_14__0
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_14__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_14__1
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_14__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM1__60_carry__1_i_14__2
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[7]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_15
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM1__60_carry__1_i_15_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_15__0
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM1__60_carry__1_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_15__1
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM1__60_carry__1_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_15__2
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM1__60_carry__1_i_15__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_1__0
       (.I0(PSUM1__60_carry__1_i_9__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_6 ),
        .I5(ALU_DIN1[13]),
        .O(PSUM1__60_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_1__1
       (.I0(PSUM1__60_carry__1_i_9__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_6 ),
        .I5(ALU_DIN1[29]),
        .O(PSUM1__60_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_1__2
       (.I0(PSUM1__60_carry__1_i_9__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_6 ),
        .I5(ALU_DIN1[13]),
        .O(PSUM1__60_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_2
       (.I0(PSUM1__60_carry__1_i_10_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_6 ),
        .I2(ALU_DIN1[29]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_7 ),
        .I5(ALU_DIN1[28]),
        .O(PSUM1__60_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_2__0
       (.I0(PSUM1__60_carry__1_i_10__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_6 ),
        .I2(ALU_DIN1[13]),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_7 ),
        .I5(ALU_DIN1[12]),
        .O(PSUM1__60_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_2__1
       (.I0(PSUM1__60_carry__1_i_10__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_6 ),
        .I2(ALU_DIN1[29]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_7 ),
        .I5(ALU_DIN1[28]),
        .O(PSUM1__60_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM1__60_carry__1_i_2__2
       (.I0(PSUM1__60_carry__1_i_10__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_6 ),
        .I2(ALU_DIN1[13]),
        .I3(ALU_DIN2[7]),
        .I4(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_7 ),
        .I5(ALU_DIN1[12]),
        .O(PSUM1__60_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM1__60_carry__1_i_3
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[29]),
        .I2(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_7 ),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[23]),
        .I5(PSUM1__60_carry__1_i_11_n_0),
        .O(PSUM1__60_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM1__60_carry__1_i_3__0
       (.I0(ALU_DIN2[22]),
        .I1(ALU_DIN1[13]),
        .I2(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_7 ),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[23]),
        .I5(PSUM1__60_carry__1_i_11__0_n_0),
        .O(PSUM1__60_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM1__60_carry__1_i_3__1
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[29]),
        .I2(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_7 ),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[7]),
        .I5(PSUM1__60_carry__1_i_11__1_n_0),
        .O(PSUM1__60_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM1__60_carry__1_i_3__2
       (.I0(ALU_DIN2[6]),
        .I1(ALU_DIN1[13]),
        .I2(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_7 ),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[7]),
        .I5(PSUM1__60_carry__1_i_11__2_n_0),
        .O(PSUM1__60_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__1_i_4
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM1__60_carry__0_i_12_n_0),
        .I5(PSUM1__60_carry__0_i_13_n_0),
        .O(PSUM1__60_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__1_i_4__0
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[22]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM1__60_carry__0_i_12__0_n_0),
        .I5(PSUM1__60_carry__0_i_13__0_n_0),
        .O(PSUM1__60_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__1_i_4__1
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM1__60_carry__0_i_12__1_n_0),
        .I5(PSUM1__60_carry__0_i_13__1_n_0),
        .O(PSUM1__60_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM1__60_carry__1_i_4__2
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[6]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM1__60_carry__0_i_12__2_n_0),
        .I5(PSUM1__60_carry__0_i_13__2_n_0),
        .O(PSUM1__60_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM1__60_carry__1_i_5
       (.I0(PSUM1__60_carry__1_i_12_n_0),
        .I1(ALU_DIN2[22]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[30]),
        .I5(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_5_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM1__60_carry__1_i_5__0
       (.I0(PSUM1__60_carry__1_i_12__0_n_0),
        .I1(ALU_DIN2[22]),
        .I2(ALU_DIN1[15]),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[14]),
        .I5(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM1__60_carry__1_i_5__1
       (.I0(PSUM1__60_carry__1_i_12__1_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[31]),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[30]),
        .I5(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM1__60_carry__1_i_5__2
       (.I0(PSUM1__60_carry__1_i_12__2_n_0),
        .I1(ALU_DIN2[6]),
        .I2(ALU_DIN1[15]),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[14]),
        .I5(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_1 ),
        .O(PSUM1__60_carry__1_i_5__2_n_0));
  LUT5 #(
    .INIT(32'h69999666)) 
    PSUM1__60_carry__1_i_6
       (.I0(PSUM1__60_carry__1_i_2_n_0),
        .I1(PSUM1__60_carry__1_i_13_n_0),
        .I2(ALU_DIN2[22]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(PSUM1__60_carry__1_i_12_n_0),
        .O(PSUM1__60_carry__1_i_6_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM1__60_carry__1_i_6__0
       (.I0(PSUM1__60_carry__1_i_2__0_n_0),
        .I1(PSUM1__60_carry__1_i_13__0_n_0),
        .I2(PSUM1__60_carry__1_i_9__0_n_0),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[13]),
        .I5(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_6__0_n_0));
  LUT5 #(
    .INIT(32'h69999666)) 
    PSUM1__60_carry__1_i_6__1
       (.I0(PSUM1__60_carry__1_i_2__1_n_0),
        .I1(PSUM1__60_carry__1_i_13__1_n_0),
        .I2(ALU_DIN2[6]),
        .I3(ALU_DIN1[31]),
        .I4(PSUM1__60_carry__1_i_12__1_n_0),
        .O(PSUM1__60_carry__1_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM1__60_carry__1_i_6__2
       (.I0(PSUM1__60_carry__1_i_2__2_n_0),
        .I1(PSUM1__60_carry__1_i_13__2_n_0),
        .I2(PSUM1__60_carry__1_i_9__2_n_0),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[13]),
        .I5(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_6 ),
        .O(PSUM1__60_carry__1_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM1__60_carry__1_i_7
       (.I0(PSUM1__60_carry__1_i_3_n_0),
        .I1(PSUM1__60_carry__1_i_14_n_0),
        .I2(PSUM1__60_carry__1_i_10_n_0),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[28]),
        .I5(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_7 ),
        .O(PSUM1__60_carry__1_i_7_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM1__60_carry__1_i_7__0
       (.I0(PSUM1__60_carry__1_i_3__0_n_0),
        .I1(PSUM1__60_carry__1_i_14__0_n_0),
        .I2(PSUM1__60_carry__1_i_10__0_n_0),
        .I3(ALU_DIN2[23]),
        .I4(ALU_DIN1[12]),
        .I5(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_7 ),
        .O(PSUM1__60_carry__1_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM1__60_carry__1_i_7__1
       (.I0(PSUM1__60_carry__1_i_3__1_n_0),
        .I1(PSUM1__60_carry__1_i_14__1_n_0),
        .I2(PSUM1__60_carry__1_i_10__1_n_0),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[28]),
        .I5(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_7 ),
        .O(PSUM1__60_carry__1_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM1__60_carry__1_i_7__2
       (.I0(PSUM1__60_carry__1_i_3__2_n_0),
        .I1(PSUM1__60_carry__1_i_14__2_n_0),
        .I2(PSUM1__60_carry__1_i_10__2_n_0),
        .I3(ALU_DIN2[7]),
        .I4(ALU_DIN1[12]),
        .I5(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_7 ),
        .O(PSUM1__60_carry__1_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM1__60_carry__1_i_8
       (.I0(PSUM1__60_carry__1_i_4_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_7 ),
        .I2(ALU_DIN1[28]),
        .I3(ALU_DIN2[23]),
        .I4(PSUM1__60_carry__1_i_15_n_0),
        .I5(PSUM1__60_carry__1_i_11_n_0),
        .O(PSUM1__60_carry__1_i_8_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM1__60_carry__1_i_8__0
       (.I0(PSUM1__60_carry__1_i_4__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_7 ),
        .I2(ALU_DIN1[12]),
        .I3(ALU_DIN2[23]),
        .I4(PSUM1__60_carry__1_i_15__0_n_0),
        .I5(PSUM1__60_carry__1_i_11__0_n_0),
        .O(PSUM1__60_carry__1_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM1__60_carry__1_i_8__1
       (.I0(PSUM1__60_carry__1_i_4__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_7 ),
        .I2(ALU_DIN1[28]),
        .I3(ALU_DIN2[7]),
        .I4(PSUM1__60_carry__1_i_15__1_n_0),
        .I5(PSUM1__60_carry__1_i_11__1_n_0),
        .O(PSUM1__60_carry__1_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM1__60_carry__1_i_8__2
       (.I0(PSUM1__60_carry__1_i_4__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_7 ),
        .I2(ALU_DIN1[12]),
        .I3(ALU_DIN2[7]),
        .I4(PSUM1__60_carry__1_i_15__2_n_0),
        .I5(PSUM1__60_carry__1_i_11__2_n_0),
        .O(PSUM1__60_carry__1_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_9
       (.I0(EX_RF_RD1[31]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[157]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM1__60_carry__1_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_9__0
       (.I0(EX_RF_RD1[15]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[141]),
        .I3(EX_RF_RD2[22]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[101]),
        .O(PSUM1__60_carry__1_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_9__1
       (.I0(EX_RF_RD1[31]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[157]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM1__60_carry__1_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM1__60_carry__1_i_9__2
       (.I0(EX_RF_RD1[15]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[141]),
        .I3(EX_RF_RD2[6]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[85]),
        .O(PSUM1__60_carry__1_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM1__60_carry__2_i_1
       (.I0(PSUM3__0_carry__0_i_10__2_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM1__60_carry__2_i_1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM1__60_carry__2_i_1__0
       (.I0(ALU_DIN1[15]),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(EX_RF_RD2[23]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[102]),
        .O(PSUM1__60_carry__2_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM1__60_carry__2_i_1__1
       (.I0(ALU_DIN1[31]),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM1__60_carry__2_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM1__60_carry__2_i_1__2
       (.I0(ALU_DIN1[15]),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(EX_RF_RD2[7]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[86]),
        .O(PSUM1__60_carry__2_i_1__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_1
       (.I0(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ),
        .O(PSUM1__60_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_1__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ),
        .O(PSUM1__60_carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_1__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ),
        .O(PSUM1__60_carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_1__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ),
        .O(PSUM1__60_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM1__60_carry_i_2
       (.I0(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ),
        .I2(ID_EX_Q[101]),
        .I3(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I4(EX_RF_RD2[22]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__60_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM1__60_carry_i_2__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ),
        .I2(ID_EX_Q[101]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[22]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__60_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM1__60_carry_i_2__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ),
        .I2(ID_EX_Q[85]),
        .I3(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I4(EX_RF_RD2[6]),
        .I5(ALU_DIN1[24]),
        .O(PSUM1__60_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM1__60_carry_i_2__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ),
        .I2(ID_EX_Q[85]),
        .I3(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I4(EX_RF_RD2[6]),
        .I5(ALU_DIN1[8]),
        .O(PSUM1__60_carry_i_2__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_3
       (.I0(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_5 ),
        .O(PSUM1__60_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_3__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_5 ),
        .O(PSUM1__60_carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_3__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_5 ),
        .O(PSUM1__60_carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_3__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_5 ),
        .O(PSUM1__60_carry_i_3__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_6 ),
        .O(PSUM1__60_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_6 ),
        .O(PSUM1__60_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_6 ),
        .O(PSUM1__60_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_6 ),
        .O(PSUM1__60_carry_i_4__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_5
       (.I0(\custom_alu/mult/mult16_3/PSUM1__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_7 ),
        .O(PSUM1__60_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_5__0
       (.I0(\custom_alu/mult/mult16_2/PSUM1__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_7 ),
        .O(PSUM1__60_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_5__1
       (.I0(\custom_alu/mult/mult16_1/PSUM1__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_7 ),
        .O(PSUM1__60_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM1__60_carry_i_5__2
       (.I0(\custom_alu/mult/mult16_0/PSUM1__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_7 ),
        .O(PSUM1__60_carry_i_5__2_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_1
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[11]),
        .O(ALU_DIN2[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_10
       (.I0(ID_EX_Q[81]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[2]),
        .O(ALU_DIN2[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_11
       (.I0(ID_EX_Q[80]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[1]),
        .O(ALU_DIN2[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_12
       (.I0(ID_EX_Q[79]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[0]),
        .O(ALU_DIN2[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_2
       (.I0(ID_EX_Q[89]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[10]),
        .O(ALU_DIN2[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_3
       (.I0(ID_EX_Q[88]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[9]),
        .O(ALU_DIN2[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_4
       (.I0(ID_EX_Q[87]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[8]),
        .O(ALU_DIN2[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_5
       (.I0(ID_EX_Q[86]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[7]),
        .O(ALU_DIN2[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_6
       (.I0(ID_EX_Q[85]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[6]),
        .O(ALU_DIN2[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_7
       (.I0(ID_EX_Q[84]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[5]),
        .O(ALU_DIN2[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_8
       (.I0(ID_EX_Q[83]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[4]),
        .O(ALU_DIN2[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM1_i_9
       (.I0(ID_EX_Q[82]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[3]),
        .O(ALU_DIN2[3]));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_1
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[22]),
        .O(PSUM2__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_10
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM2__0_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_10__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM2__0_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_10__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM2__0_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_10__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM2__0_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_11
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[25]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[104]),
        .O(PSUM2__0_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_11__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[25]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[104]),
        .O(PSUM2__0_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_11__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[9]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[88]),
        .O(PSUM2__0_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_11__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[9]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[88]),
        .O(PSUM2__0_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_12
       (.I0(EX_RF_RD1[18]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[144]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM2__0_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_12__0
       (.I0(EX_RF_RD1[2]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[128]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM2__0_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_12__1
       (.I0(EX_RF_RD1[18]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[144]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM2__0_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_12__2
       (.I0(EX_RF_RD1[2]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[128]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM2__0_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_1__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[6]),
        .O(PSUM2__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_1__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[22]),
        .O(PSUM2__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_1__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[6]),
        .O(PSUM2__0_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_2
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[21]),
        .O(PSUM2__0_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_2__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[5]),
        .O(PSUM2__0_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_2__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[21]),
        .O(PSUM2__0_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_2__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[5]),
        .O(PSUM2__0_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_3
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[20]),
        .O(PSUM2__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_3__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[4]),
        .O(PSUM2__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_3__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[20]),
        .O(PSUM2__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_3__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[4]),
        .O(PSUM2__0_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_4
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[19]),
        .O(PSUM2__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_4__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[3]),
        .O(PSUM2__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_4__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[19]),
        .O(PSUM2__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__0_i_4__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[3]),
        .O(PSUM2__0_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_5
       (.I0(PSUM2__0_carry__0_i_1_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM2__0_carry__0_i_9_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_5__0
       (.I0(PSUM2__0_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM2__0_carry__0_i_9__0_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_5__1
       (.I0(PSUM2__0_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM2__0_carry__0_i_9__1_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_5__2
       (.I0(PSUM2__0_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM2__0_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_6
       (.I0(PSUM2__0_carry__0_i_2_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM2__0_carry__0_i_10_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_6__0
       (.I0(PSUM2__0_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM2__0_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_6__1
       (.I0(PSUM2__0_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM2__0_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_6__2
       (.I0(PSUM2__0_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM2__0_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__0_carry__0_i_7
       (.I0(PSUM2__0_carry__0_i_3_n_0),
        .I1(PSUM2__0_carry__0_i_11_n_0),
        .I2(ALU_DIN2[26]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__0_carry__0_i_7__0
       (.I0(PSUM2__0_carry__0_i_3__0_n_0),
        .I1(PSUM2__0_carry__0_i_11__0_n_0),
        .I2(ALU_DIN2[26]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__0_carry__0_i_7__1
       (.I0(PSUM2__0_carry__0_i_3__1_n_0),
        .I1(PSUM2__0_carry__0_i_11__1_n_0),
        .I2(ALU_DIN2[10]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__0_carry__0_i_7__2
       (.I0(PSUM2__0_carry__0_i_3__2_n_0),
        .I1(PSUM2__0_carry__0_i_11__2_n_0),
        .I2(ALU_DIN2[10]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_8
       (.I0(PSUM2__0_carry__0_i_4_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[19]),
        .I3(PSUM2__0_carry__0_i_12_n_0),
        .I4(ALU_DIN1[20]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_8__0
       (.I0(PSUM2__0_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[3]),
        .I3(PSUM2__0_carry__0_i_12__0_n_0),
        .I4(ALU_DIN1[4]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_8__1
       (.I0(PSUM2__0_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[19]),
        .I3(PSUM2__0_carry__0_i_12__1_n_0),
        .I4(ALU_DIN1[20]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__0_carry__0_i_8__2
       (.I0(PSUM2__0_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[3]),
        .I3(PSUM2__0_carry__0_i_12__2_n_0),
        .I4(ALU_DIN1[4]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_9
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM2__0_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_9__0
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM2__0_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_9__1
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM2__0_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry__0_i_9__2
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM2__0_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__0_carry__1_i_1
       (.I0(ID_EX_Q[105]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[26]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[25]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__0_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__0_carry__1_i_1__0
       (.I0(ID_EX_Q[105]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[26]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[25]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__0_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__0_carry__1_i_1__1
       (.I0(ID_EX_Q[89]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[10]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[9]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__0_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__0_carry__1_i_1__2
       (.I0(ID_EX_Q[89]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[10]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[9]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__0_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__1_i_2
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__0_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__1_i_2__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__0_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__1_i_2__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__0_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__0_carry__1_i_2__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__0_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__0_carry__1_i_3
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__0_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__0_carry__1_i_3__0
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__0_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__0_carry__1_i_3__1
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[88]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[10]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__0_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__0_carry__1_i_3__2
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[88]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[10]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__0_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__0_carry__1_i_4
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[26]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[25]),
        .O(PSUM2__0_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__0_carry__1_i_4__0
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[26]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[25]),
        .O(PSUM2__0_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__0_carry__1_i_4__1
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[10]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[9]),
        .O(PSUM2__0_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__0_carry__1_i_4__2
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[10]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[9]),
        .O(PSUM2__0_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_1
       (.I0(ALU_DIN2[25]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[26]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_1__0
       (.I0(ALU_DIN2[25]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[26]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[24]),
        .O(PSUM2__0_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_1__1
       (.I0(ALU_DIN2[9]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[10]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_1__2
       (.I0(ALU_DIN2[9]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[10]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[8]),
        .O(PSUM2__0_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__0_carry_i_2
       (.I0(ID_EX_Q[104]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[25]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__0_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__0_carry_i_2__0
       (.I0(ID_EX_Q[104]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[25]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__0_carry_i_2__1
       (.I0(ID_EX_Q[88]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[9]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[10]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__0_carry_i_2__2
       (.I0(ID_EX_Q[88]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[9]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[10]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__0_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__0_carry_i_3
       (.I0(ID_EX_Q[103]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[24]),
        .I3(ID_EX_Q[143]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[17]),
        .O(PSUM2__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__0_carry_i_3__0
       (.I0(ID_EX_Q[103]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[24]),
        .I3(ID_EX_Q[127]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[1]),
        .O(PSUM2__0_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__0_carry_i_3__1
       (.I0(ID_EX_Q[87]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[8]),
        .I3(ID_EX_Q[143]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[17]),
        .O(PSUM2__0_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__0_carry_i_3__2
       (.I0(ID_EX_Q[87]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[8]),
        .I3(ID_EX_Q[127]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[1]),
        .O(PSUM2__0_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__0_carry_i_4
       (.I0(ALU_DIN1[18]),
        .I1(PSUM2__0_carry_i_8_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[26]),
        .O(PSUM2__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__0_carry_i_4__0
       (.I0(ALU_DIN1[2]),
        .I1(PSUM2__0_carry_i_8__0_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[26]),
        .O(PSUM2__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__0_carry_i_4__1
       (.I0(ALU_DIN1[18]),
        .I1(PSUM2__0_carry_i_8__1_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[10]),
        .O(PSUM2__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__0_carry_i_4__2
       (.I0(ALU_DIN1[2]),
        .I1(PSUM2__0_carry_i_8__2_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[10]),
        .O(PSUM2__0_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_5
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[26]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[18]),
        .O(PSUM2__0_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_5__0
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[26]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[2]),
        .O(PSUM2__0_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_5__1
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[10]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[18]),
        .O(PSUM2__0_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__0_carry_i_5__2
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[10]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[2]),
        .O(PSUM2__0_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM2__0_carry_i_6
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[17]),
        .I2(ID_EX_Q[104]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[25]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__0_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM2__0_carry_i_6__0
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[1]),
        .I2(ID_EX_Q[104]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[25]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__0_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM2__0_carry_i_6__1
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[17]),
        .I2(ID_EX_Q[88]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[9]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__0_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM2__0_carry_i_6__2
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[1]),
        .I2(ID_EX_Q[88]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[9]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__0_carry_i_6__2_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__0_carry_i_7
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM2__0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__0_carry_i_7__0
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM2__0_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__0_carry_i_7__1
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM2__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__0_carry_i_7__2
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM2__0_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry_i_8
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM2__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry_i_8__0
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM2__0_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry_i_8__1
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM2__0_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__0_carry_i_8__2
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM2__0_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_1
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[22]),
        .O(PSUM2__30_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_10
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM2__30_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_10__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM2__30_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_10__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM2__30_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_10__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM2__30_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_11
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[28]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[107]),
        .O(PSUM2__30_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_11__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[28]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[107]),
        .O(PSUM2__30_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_11__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[12]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[91]),
        .O(PSUM2__30_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_11__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[12]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[91]),
        .O(PSUM2__30_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_12
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM2__30_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_12__0
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM2__30_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_12__1
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[146]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM2__30_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_12__2
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM2__30_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_1__0
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[6]),
        .O(PSUM2__30_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_1__1
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[20]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[22]),
        .O(PSUM2__30_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_1__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[4]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[5]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[6]),
        .O(PSUM2__30_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_2
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[21]),
        .O(PSUM2__30_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_2__0
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[5]),
        .O(PSUM2__30_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_2__1
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[19]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[21]),
        .O(PSUM2__30_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_2__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[5]),
        .O(PSUM2__30_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_3
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[20]),
        .O(PSUM2__30_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_3__0
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[4]),
        .O(PSUM2__30_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_3__1
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[20]),
        .O(PSUM2__30_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_3__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[4]),
        .O(PSUM2__30_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_4
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[19]),
        .O(PSUM2__30_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_4__0
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[3]),
        .O(PSUM2__30_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_4__1
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[19]),
        .O(PSUM2__30_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__0_i_4__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[3]),
        .O(PSUM2__30_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_5
       (.I0(PSUM2__30_carry__0_i_1_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM2__30_carry__0_i_9_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_5__0
       (.I0(PSUM2__30_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM2__30_carry__0_i_9__0_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_5__1
       (.I0(PSUM2__30_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM2__30_carry__0_i_9__1_n_0),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_5__2
       (.I0(PSUM2__30_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[6]),
        .I3(PSUM2__30_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_6
       (.I0(PSUM2__30_carry__0_i_2_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM2__30_carry__0_i_10_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_6__0
       (.I0(PSUM2__30_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM2__30_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_6__1
       (.I0(PSUM2__30_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[21]),
        .I3(PSUM2__30_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM2__30_carry__0_i_6__2
       (.I0(PSUM2__30_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[5]),
        .I3(PSUM2__30_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__30_carry__0_i_7
       (.I0(PSUM2__30_carry__0_i_3_n_0),
        .I1(PSUM2__30_carry__0_i_11_n_0),
        .I2(ALU_DIN2[29]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__30_carry__0_i_7__0
       (.I0(PSUM2__30_carry__0_i_3__0_n_0),
        .I1(PSUM2__30_carry__0_i_11__0_n_0),
        .I2(ALU_DIN2[29]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__30_carry__0_i_7__1
       (.I0(PSUM2__30_carry__0_i_3__1_n_0),
        .I1(PSUM2__30_carry__0_i_11__1_n_0),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN1[19]),
        .I4(ALU_DIN1[21]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM2__30_carry__0_i_7__2
       (.I0(PSUM2__30_carry__0_i_3__2_n_0),
        .I1(PSUM2__30_carry__0_i_11__2_n_0),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN1[3]),
        .I4(ALU_DIN1[5]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A6A6A959595)) 
    PSUM2__30_carry__0_i_8
       (.I0(PSUM2__30_carry__0_i_4_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[19]),
        .I3(ALU_DIN2[29]),
        .I4(ALU_DIN1[18]),
        .I5(PSUM2__30_carry__0_i_12_n_0),
        .O(PSUM2__30_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A6A6A959595)) 
    PSUM2__30_carry__0_i_8__0
       (.I0(PSUM2__30_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[3]),
        .I3(ALU_DIN2[29]),
        .I4(ALU_DIN1[2]),
        .I5(PSUM2__30_carry__0_i_12__0_n_0),
        .O(PSUM2__30_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A6A6A959595)) 
    PSUM2__30_carry__0_i_8__1
       (.I0(PSUM2__30_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[19]),
        .I3(ALU_DIN2[13]),
        .I4(ALU_DIN1[18]),
        .I5(PSUM2__30_carry__0_i_12__1_n_0),
        .O(PSUM2__30_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A6A6A959595)) 
    PSUM2__30_carry__0_i_8__2
       (.I0(PSUM2__30_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[3]),
        .I3(ALU_DIN2[13]),
        .I4(ALU_DIN1[2]),
        .I5(PSUM2__30_carry__0_i_12__2_n_0),
        .O(PSUM2__30_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_9
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM2__30_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_9__0
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM2__30_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_9__1
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM2__30_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry__0_i_9__2
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM2__30_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__30_carry__1_i_1
       (.I0(ID_EX_Q[108]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[29]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__30_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__30_carry__1_i_1__0
       (.I0(ID_EX_Q[108]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[29]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__30_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__30_carry__1_i_1__1
       (.I0(ID_EX_Q[92]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[13]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[12]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__30_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM2__30_carry__1_i_1__2
       (.I0(ID_EX_Q[92]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[13]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[12]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__30_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__1_i_2
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__30_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__1_i_2__0
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__30_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__1_i_2__1
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__30_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM2__30_carry__1_i_2__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__30_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__30_carry__1_i_3
       (.I0(EX_RF_RD2[28]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[107]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[29]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__30_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__30_carry__1_i_3__0
       (.I0(EX_RF_RD2[28]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[107]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[29]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__30_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__30_carry__1_i_3__1
       (.I0(EX_RF_RD2[12]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[91]),
        .I3(ALU_DIN1[22]),
        .I4(ALU_DIN2[13]),
        .I5(ALU_DIN1[23]),
        .O(PSUM2__30_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM2__30_carry__1_i_3__2
       (.I0(EX_RF_RD2[12]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[91]),
        .I3(ALU_DIN1[6]),
        .I4(ALU_DIN2[13]),
        .I5(ALU_DIN1[7]),
        .O(PSUM2__30_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__30_carry__1_i_4
       (.I0(ALU_DIN2[27]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[29]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[28]),
        .O(PSUM2__30_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__30_carry__1_i_4__0
       (.I0(ALU_DIN2[27]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[29]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[28]),
        .O(PSUM2__30_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__30_carry__1_i_4__1
       (.I0(ALU_DIN2[11]),
        .I1(ALU_DIN1[21]),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[13]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN2[12]),
        .O(PSUM2__30_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM2__30_carry__1_i_4__2
       (.I0(ALU_DIN2[11]),
        .I1(ALU_DIN1[5]),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[13]),
        .I4(ALU_DIN1[7]),
        .I5(ALU_DIN2[12]),
        .O(PSUM2__30_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_1
       (.I0(ALU_DIN2[28]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[29]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_1__0
       (.I0(ALU_DIN2[28]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[29]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[27]),
        .O(PSUM2__30_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_1__1
       (.I0(ALU_DIN2[12]),
        .I1(ALU_DIN1[18]),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN1[19]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_1__2
       (.I0(ALU_DIN2[12]),
        .I1(ALU_DIN1[2]),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN2[11]),
        .O(PSUM2__30_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_2
       (.I0(ID_EX_Q[107]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[28]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[29]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__30_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_2__0
       (.I0(ID_EX_Q[107]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[28]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[29]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__30_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_2__1
       (.I0(ID_EX_Q[91]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[12]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[13]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__30_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_2__2
       (.I0(ID_EX_Q[91]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[12]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[13]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__30_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__30_carry_i_3
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ID_EX_Q[143]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[17]),
        .O(PSUM2__30_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__30_carry_i_3__0
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ID_EX_Q[127]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[1]),
        .O(PSUM2__30_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__30_carry_i_3__1
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ID_EX_Q[143]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[17]),
        .O(PSUM2__30_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM2__30_carry_i_3__2
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ID_EX_Q[127]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[1]),
        .O(PSUM2__30_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__30_carry_i_4
       (.I0(ALU_DIN1[18]),
        .I1(PSUM2__30_carry_i_8_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[29]),
        .O(PSUM2__30_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__30_carry_i_4__0
       (.I0(ALU_DIN1[2]),
        .I1(PSUM2__30_carry_i_8__0_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[29]),
        .O(PSUM2__30_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__30_carry_i_4__1
       (.I0(ALU_DIN1[18]),
        .I1(PSUM2__30_carry_i_8__1_n_0),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[13]),
        .O(PSUM2__30_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM2__30_carry_i_4__2
       (.I0(ALU_DIN1[2]),
        .I1(PSUM2__30_carry_i_8__2_n_0),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[13]),
        .O(PSUM2__30_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_5
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[29]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[18]),
        .O(PSUM2__30_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_5__0
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[29]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[2]),
        .O(PSUM2__30_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_5__1
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[13]),
        .I2(ALU_DIN1[17]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[18]),
        .O(PSUM2__30_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM2__30_carry_i_5__2
       (.I0(ALU_DIN1[0]),
        .I1(ALU_DIN2[13]),
        .I2(ALU_DIN1[1]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[2]),
        .O(PSUM2__30_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_6
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__30_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_6__0
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__30_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_6__1
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[12]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__30_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM2__30_carry_i_6__2
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ALU_DIN1[1]),
        .I4(ALU_DIN2[12]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__30_carry_i_6__2_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__30_carry_i_7
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM2__30_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__30_carry_i_7__0
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM2__30_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__30_carry_i_7__1
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM2__30_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM2__30_carry_i_7__2
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM2__30_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry_i_8
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM2__30_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry_i_8__0
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM2__30_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry_i_8__1
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM2__30_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__30_carry_i_8__2
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[129]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM2__30_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__0_i_1
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM2__60_carry__0_i_9_n_0),
        .I5(PSUM2__60_carry__0_i_10_n_0),
        .O(PSUM2__60_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_10
       (.I0(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_7 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[17]),
        .O(PSUM2__60_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_10__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_7 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[1]),
        .O(PSUM2__60_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_10__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_7 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[17]),
        .O(PSUM2__60_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_10__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_7 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[1]),
        .O(PSUM2__60_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_11
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_7 ),
        .O(PSUM2__60_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_11__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_7 ),
        .O(PSUM2__60_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_11__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_7 ),
        .O(PSUM2__60_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_11__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_7 ),
        .O(PSUM2__60_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_12
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[19]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_1 ),
        .O(PSUM2__60_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_12__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[3]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_1 ),
        .O(PSUM2__60_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_12__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[19]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_1 ),
        .O(PSUM2__60_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_12__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[3]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_1 ),
        .O(PSUM2__60_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_13
       (.I0(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_6 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[18]),
        .O(PSUM2__60_carry__0_i_13_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_13__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_6 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[2]),
        .O(PSUM2__60_carry__0_i_13__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_13__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_6 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[18]),
        .O(PSUM2__60_carry__0_i_13__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__0_i_13__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_6 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[2]),
        .O(PSUM2__60_carry__0_i_13__2_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM2__60_carry__0_i_14
       (.I0(ALU_DIN1[17]),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[30]),
        .I5(PSUM2__60_carry__0_i_11_n_0),
        .O(PSUM2__60_carry__0_i_14_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM2__60_carry__0_i_14__0
       (.I0(ALU_DIN1[1]),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[30]),
        .I5(PSUM2__60_carry__0_i_11__0_n_0),
        .O(PSUM2__60_carry__0_i_14__0_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM2__60_carry__0_i_14__1
       (.I0(ALU_DIN1[17]),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ),
        .I3(ALU_DIN1[18]),
        .I4(ALU_DIN2[14]),
        .I5(PSUM2__60_carry__0_i_11__1_n_0),
        .O(PSUM2__60_carry__0_i_14__1_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM2__60_carry__0_i_14__2
       (.I0(ALU_DIN1[1]),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ),
        .I3(ALU_DIN1[2]),
        .I4(ALU_DIN2[14]),
        .I5(PSUM2__60_carry__0_i_11__2_n_0),
        .O(PSUM2__60_carry__0_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_15
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[16]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_4 ),
        .O(PSUM2__60_carry__0_i_15_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_15__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[0]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_4 ),
        .O(PSUM2__60_carry__0_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_15__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[16]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_4 ),
        .O(PSUM2__60_carry__0_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_15__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[0]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_4 ),
        .O(PSUM2__60_carry__0_i_15__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__0_i_1__0
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM2__60_carry__0_i_9__0_n_0),
        .I5(PSUM2__60_carry__0_i_10__0_n_0),
        .O(PSUM2__60_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__0_i_1__1
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM2__60_carry__0_i_9__1_n_0),
        .I5(PSUM2__60_carry__0_i_10__1_n_0),
        .O(PSUM2__60_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__0_i_1__2
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM2__60_carry__0_i_9__2_n_0),
        .I5(PSUM2__60_carry__0_i_10__2_n_0),
        .O(PSUM2__60_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM2__60_carry__0_i_2
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[18]),
        .I2(PSUM2__60_carry__0_i_11_n_0),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM2__60_carry__0_i_2__0
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[2]),
        .I2(PSUM2__60_carry__0_i_11__0_n_0),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM2__60_carry__0_i_2__1
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[18]),
        .I2(PSUM2__60_carry__0_i_11__1_n_0),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM2__60_carry__0_i_2__2
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[2]),
        .I2(PSUM2__60_carry__0_i_11__2_n_0),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM2__60_carry__0_i_3
       (.I0(PSUM2__60_carry__0_i_11_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN1[18]),
        .I3(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ),
        .I5(ALU_DIN1[17]),
        .O(PSUM2__60_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM2__60_carry__0_i_3__0
       (.I0(PSUM2__60_carry__0_i_11__0_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN1[2]),
        .I3(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ),
        .I5(ALU_DIN1[1]),
        .O(PSUM2__60_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM2__60_carry__0_i_3__1
       (.I0(PSUM2__60_carry__0_i_11__1_n_0),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN1[18]),
        .I3(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ),
        .I5(ALU_DIN1[17]),
        .O(PSUM2__60_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM2__60_carry__0_i_3__2
       (.I0(PSUM2__60_carry__0_i_11__2_n_0),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN1[2]),
        .I3(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ),
        .I5(ALU_DIN1[1]),
        .O(PSUM2__60_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM2__60_carry__0_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_7 ),
        .I2(ALU_DIN1[16]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM2__60_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM2__60_carry__0_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_7 ),
        .I2(ALU_DIN1[0]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM2__60_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM2__60_carry__0_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_7 ),
        .I2(ALU_DIN1[16]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM2__60_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM2__60_carry__0_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_7 ),
        .I2(ALU_DIN1[0]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM2__60_carry__0_i_4__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_5
       (.I0(PSUM2__60_carry__0_i_1_n_0),
        .I1(PSUM2__60_carry__0_i_12_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM2__60_carry__0_i_13_n_0),
        .O(PSUM2__60_carry__0_i_5_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_5__0
       (.I0(PSUM2__60_carry__0_i_1__0_n_0),
        .I1(PSUM2__60_carry__0_i_12__0_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM2__60_carry__0_i_13__0_n_0),
        .O(PSUM2__60_carry__0_i_5__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_5__1
       (.I0(PSUM2__60_carry__0_i_1__1_n_0),
        .I1(PSUM2__60_carry__0_i_12__1_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM2__60_carry__0_i_13__1_n_0),
        .O(PSUM2__60_carry__0_i_5__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_5__2
       (.I0(PSUM2__60_carry__0_i_1__2_n_0),
        .I1(PSUM2__60_carry__0_i_12__2_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM2__60_carry__0_i_13__2_n_0),
        .O(PSUM2__60_carry__0_i_5__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_6
       (.I0(PSUM2__60_carry__0_i_2_n_0),
        .I1(PSUM2__60_carry__0_i_9_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM2__60_carry__0_i_10_n_0),
        .O(PSUM2__60_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_6__0
       (.I0(PSUM2__60_carry__0_i_2__0_n_0),
        .I1(PSUM2__60_carry__0_i_9__0_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM2__60_carry__0_i_10__0_n_0),
        .O(PSUM2__60_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_6__1
       (.I0(PSUM2__60_carry__0_i_2__1_n_0),
        .I1(PSUM2__60_carry__0_i_9__1_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[19]),
        .I4(PSUM2__60_carry__0_i_10__1_n_0),
        .O(PSUM2__60_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM2__60_carry__0_i_6__2
       (.I0(PSUM2__60_carry__0_i_2__2_n_0),
        .I1(PSUM2__60_carry__0_i_9__2_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[3]),
        .I4(PSUM2__60_carry__0_i_10__2_n_0),
        .O(PSUM2__60_carry__0_i_6__2_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM2__60_carry__0_i_7
       (.I0(PSUM2__60_carry__0_i_14_n_0),
        .I1(ALU_DIN1[16]),
        .I2(ALU_DIN2[31]),
        .I3(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_7 ),
        .O(PSUM2__60_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM2__60_carry__0_i_7__0
       (.I0(PSUM2__60_carry__0_i_14__0_n_0),
        .I1(ALU_DIN1[0]),
        .I2(ALU_DIN2[31]),
        .I3(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_7 ),
        .O(PSUM2__60_carry__0_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM2__60_carry__0_i_7__1
       (.I0(PSUM2__60_carry__0_i_14__1_n_0),
        .I1(ALU_DIN1[16]),
        .I2(ALU_DIN2[15]),
        .I3(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_7 ),
        .O(PSUM2__60_carry__0_i_7__1_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM2__60_carry__0_i_7__2
       (.I0(PSUM2__60_carry__0_i_14__2_n_0),
        .I1(ALU_DIN1[0]),
        .I2(ALU_DIN2[15]),
        .I3(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_7 ),
        .O(PSUM2__60_carry__0_i_7__2_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM2__60_carry__0_i_8
       (.I0(PSUM2__60_carry__0_i_15_n_0),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[30]),
        .I3(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_8_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM2__60_carry__0_i_8__0
       (.I0(PSUM2__60_carry__0_i_15__0_n_0),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[30]),
        .I3(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM2__60_carry__0_i_8__1
       (.I0(PSUM2__60_carry__0_i_15__1_n_0),
        .I1(ALU_DIN1[17]),
        .I2(ALU_DIN2[14]),
        .I3(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM2__60_carry__0_i_8__2
       (.I0(PSUM2__60_carry__0_i_15__2_n_0),
        .I1(ALU_DIN1[1]),
        .I2(ALU_DIN2[14]),
        .I3(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ),
        .O(PSUM2__60_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_9
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[18]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_6 ),
        .O(PSUM2__60_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_9__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[2]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_6 ),
        .O(PSUM2__60_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_9__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[18]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_6 ),
        .O(PSUM2__60_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM2__60_carry__0_i_9__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[2]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_6 ),
        .O(PSUM2__60_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_1
       (.I0(PSUM2__60_carry__1_i_9_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_6 ),
        .I5(ALU_DIN1[21]),
        .O(PSUM2__60_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_10
       (.I0(EX_RF_RD1[22]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[148]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM2__60_carry__1_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_10__0
       (.I0(EX_RF_RD1[6]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[132]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM2__60_carry__1_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_10__1
       (.I0(EX_RF_RD1[22]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[148]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM2__60_carry__1_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_10__2
       (.I0(EX_RF_RD1[6]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[132]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM2__60_carry__1_i_10__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__1_i_11
       (.I0(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_1 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[19]),
        .O(PSUM2__60_carry__1_i_11_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__1_i_11__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_1 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[3]),
        .O(PSUM2__60_carry__1_i_11__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__1_i_11__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_1 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[19]),
        .O(PSUM2__60_carry__1_i_11__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM2__60_carry__1_i_11__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_1 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[3]),
        .O(PSUM2__60_carry__1_i_11__2_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_12
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[21]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_6 ),
        .O(PSUM2__60_carry__1_i_12_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_12__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[5]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_6 ),
        .O(PSUM2__60_carry__1_i_12__0_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_12__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[21]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_6 ),
        .O(PSUM2__60_carry__1_i_12__1_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_12__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[5]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_6 ),
        .O(PSUM2__60_carry__1_i_12__2_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM2__60_carry__1_i_13
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[22]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM2__60_carry__1_i_13__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[6]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_13__0_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM2__60_carry__1_i_13__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[22]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_13__1_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM2__60_carry__1_i_13__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[6]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_13__2_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_14
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[20]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_7 ),
        .O(PSUM2__60_carry__1_i_14_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_14__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[4]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_7 ),
        .O(PSUM2__60_carry__1_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_14__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[20]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_7 ),
        .O(PSUM2__60_carry__1_i_14__1_n_0));
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM2__60_carry__1_i_14__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[4]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_7 ),
        .O(PSUM2__60_carry__1_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_15
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM2__60_carry__1_i_15_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_15__0
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM2__60_carry__1_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_15__1
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[147]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM2__60_carry__1_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_15__2
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM2__60_carry__1_i_15__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_1__0
       (.I0(PSUM2__60_carry__1_i_9__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_6 ),
        .I5(ALU_DIN1[5]),
        .O(PSUM2__60_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_1__1
       (.I0(PSUM2__60_carry__1_i_9__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_6 ),
        .I5(ALU_DIN1[21]),
        .O(PSUM2__60_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_1__2
       (.I0(PSUM2__60_carry__1_i_9__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_6 ),
        .I5(ALU_DIN1[5]),
        .O(PSUM2__60_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_2
       (.I0(PSUM2__60_carry__1_i_10_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_7 ),
        .I5(ALU_DIN1[20]),
        .O(PSUM2__60_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_2__0
       (.I0(PSUM2__60_carry__1_i_10__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_7 ),
        .I5(ALU_DIN1[4]),
        .O(PSUM2__60_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_2__1
       (.I0(PSUM2__60_carry__1_i_10__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_7 ),
        .I5(ALU_DIN1[20]),
        .O(PSUM2__60_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM2__60_carry__1_i_2__2
       (.I0(PSUM2__60_carry__1_i_10__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_7 ),
        .I5(ALU_DIN1[4]),
        .O(PSUM2__60_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM2__60_carry__1_i_3
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[21]),
        .I2(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_7 ),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[31]),
        .I5(PSUM2__60_carry__1_i_11_n_0),
        .O(PSUM2__60_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM2__60_carry__1_i_3__0
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[5]),
        .I2(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_7 ),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[31]),
        .I5(PSUM2__60_carry__1_i_11__0_n_0),
        .O(PSUM2__60_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM2__60_carry__1_i_3__1
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[21]),
        .I2(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_7 ),
        .I3(ALU_DIN1[20]),
        .I4(ALU_DIN2[15]),
        .I5(PSUM2__60_carry__1_i_11__1_n_0),
        .O(PSUM2__60_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM2__60_carry__1_i_3__2
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[5]),
        .I2(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_7 ),
        .I3(ALU_DIN1[4]),
        .I4(ALU_DIN2[15]),
        .I5(PSUM2__60_carry__1_i_11__2_n_0),
        .O(PSUM2__60_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__1_i_4
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM2__60_carry__0_i_12_n_0),
        .I5(PSUM2__60_carry__0_i_13_n_0),
        .O(PSUM2__60_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__1_i_4__0
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM2__60_carry__0_i_12__0_n_0),
        .I5(PSUM2__60_carry__0_i_13__0_n_0),
        .O(PSUM2__60_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__1_i_4__1
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[20]),
        .I4(PSUM2__60_carry__0_i_12__1_n_0),
        .I5(PSUM2__60_carry__0_i_13__1_n_0),
        .O(PSUM2__60_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM2__60_carry__1_i_4__2
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[4]),
        .I4(PSUM2__60_carry__0_i_12__2_n_0),
        .I5(PSUM2__60_carry__0_i_13__2_n_0),
        .O(PSUM2__60_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM2__60_carry__1_i_5
       (.I0(PSUM2__60_carry__1_i_12_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN2[31]),
        .I4(ALU_DIN1[22]),
        .I5(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_5_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM2__60_carry__1_i_5__0
       (.I0(PSUM2__60_carry__1_i_12__0_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN1[7]),
        .I3(ALU_DIN2[31]),
        .I4(ALU_DIN1[6]),
        .I5(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM2__60_carry__1_i_5__1
       (.I0(PSUM2__60_carry__1_i_12__1_n_0),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[22]),
        .I5(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM2__60_carry__1_i_5__2
       (.I0(PSUM2__60_carry__1_i_12__2_n_0),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN1[7]),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[6]),
        .I5(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_1 ),
        .O(PSUM2__60_carry__1_i_5__2_n_0));
  LUT5 #(
    .INIT(32'h69999666)) 
    PSUM2__60_carry__1_i_6
       (.I0(PSUM2__60_carry__1_i_2_n_0),
        .I1(PSUM2__60_carry__1_i_13_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[23]),
        .I4(PSUM2__60_carry__1_i_12_n_0),
        .O(PSUM2__60_carry__1_i_6_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM2__60_carry__1_i_6__0
       (.I0(PSUM2__60_carry__1_i_2__0_n_0),
        .I1(PSUM2__60_carry__1_i_13__0_n_0),
        .I2(PSUM2__60_carry__1_i_9__0_n_0),
        .I3(ALU_DIN2[31]),
        .I4(ALU_DIN1[5]),
        .I5(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_6 ),
        .O(PSUM2__60_carry__1_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM2__60_carry__1_i_6__1
       (.I0(PSUM2__60_carry__1_i_2__1_n_0),
        .I1(PSUM2__60_carry__1_i_13__1_n_0),
        .I2(PSUM2__60_carry__1_i_9__1_n_0),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[21]),
        .I5(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_6 ),
        .O(PSUM2__60_carry__1_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM2__60_carry__1_i_6__2
       (.I0(PSUM2__60_carry__1_i_2__2_n_0),
        .I1(PSUM2__60_carry__1_i_13__2_n_0),
        .I2(PSUM2__60_carry__1_i_9__2_n_0),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[5]),
        .I5(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_6 ),
        .O(PSUM2__60_carry__1_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM2__60_carry__1_i_7
       (.I0(PSUM2__60_carry__1_i_3_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[31]),
        .I4(PSUM2__60_carry__1_i_10_n_0),
        .I5(PSUM2__60_carry__1_i_14_n_0),
        .O(PSUM2__60_carry__1_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM2__60_carry__1_i_7__0
       (.I0(PSUM2__60_carry__1_i_3__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[31]),
        .I4(PSUM2__60_carry__1_i_10__0_n_0),
        .I5(PSUM2__60_carry__1_i_14__0_n_0),
        .O(PSUM2__60_carry__1_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM2__60_carry__1_i_7__1
       (.I0(PSUM2__60_carry__1_i_3__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[21]),
        .I3(ALU_DIN2[15]),
        .I4(PSUM2__60_carry__1_i_10__1_n_0),
        .I5(PSUM2__60_carry__1_i_14__1_n_0),
        .O(PSUM2__60_carry__1_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h9666699969999666)) 
    PSUM2__60_carry__1_i_7__2
       (.I0(PSUM2__60_carry__1_i_3__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_6 ),
        .I2(ALU_DIN1[5]),
        .I3(ALU_DIN2[15]),
        .I4(PSUM2__60_carry__1_i_10__2_n_0),
        .I5(PSUM2__60_carry__1_i_14__2_n_0),
        .O(PSUM2__60_carry__1_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM2__60_carry__1_i_8
       (.I0(PSUM2__60_carry__1_i_4_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_7 ),
        .I2(ALU_DIN1[20]),
        .I3(ALU_DIN2[31]),
        .I4(PSUM2__60_carry__1_i_15_n_0),
        .I5(PSUM2__60_carry__1_i_11_n_0),
        .O(PSUM2__60_carry__1_i_8_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM2__60_carry__1_i_8__0
       (.I0(PSUM2__60_carry__1_i_4__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_7 ),
        .I2(ALU_DIN1[4]),
        .I3(ALU_DIN2[31]),
        .I4(PSUM2__60_carry__1_i_15__0_n_0),
        .I5(PSUM2__60_carry__1_i_11__0_n_0),
        .O(PSUM2__60_carry__1_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM2__60_carry__1_i_8__1
       (.I0(PSUM2__60_carry__1_i_4__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_7 ),
        .I2(ALU_DIN1[20]),
        .I3(ALU_DIN2[15]),
        .I4(PSUM2__60_carry__1_i_15__1_n_0),
        .I5(PSUM2__60_carry__1_i_11__1_n_0),
        .O(PSUM2__60_carry__1_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM2__60_carry__1_i_8__2
       (.I0(PSUM2__60_carry__1_i_4__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_7 ),
        .I2(ALU_DIN1[4]),
        .I3(ALU_DIN2[15]),
        .I4(PSUM2__60_carry__1_i_15__2_n_0),
        .I5(PSUM2__60_carry__1_i_11__2_n_0),
        .O(PSUM2__60_carry__1_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_9
       (.I0(EX_RF_RD1[23]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[149]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM2__60_carry__1_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_9__0
       (.I0(EX_RF_RD1[7]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[133]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM2__60_carry__1_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_9__1
       (.I0(EX_RF_RD1[23]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[149]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM2__60_carry__1_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM2__60_carry__1_i_9__2
       (.I0(EX_RF_RD1[7]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[133]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM2__60_carry__1_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM2__60_carry__2_i_1
       (.I0(ALU_DIN1[23]),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM2__60_carry__2_i_1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM2__60_carry__2_i_1__0
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM2__60_carry__2_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM2__60_carry__2_i_1__1
       (.I0(ALU_DIN1[23]),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[22]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM2__60_carry__2_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM2__60_carry__2_i_1__2
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_1 ),
        .I2(ALU_DIN1[6]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM2__60_carry__2_i_1__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_1
       (.I0(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ),
        .O(PSUM2__60_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_1__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ),
        .O(PSUM2__60_carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_1__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ),
        .O(PSUM2__60_carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_1__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ),
        .O(PSUM2__60_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM2__60_carry_i_2
       (.I0(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ),
        .I2(ID_EX_Q[109]),
        .I3(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I4(EX_RF_RD2[30]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__60_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM2__60_carry_i_2__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ),
        .I2(ID_EX_Q[109]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[30]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__60_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM2__60_carry_i_2__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ),
        .I2(ID_EX_Q[93]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[14]),
        .I5(ALU_DIN1[16]),
        .O(PSUM2__60_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM2__60_carry_i_2__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ),
        .I2(ID_EX_Q[93]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[14]),
        .I5(ALU_DIN1[0]),
        .O(PSUM2__60_carry_i_2__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_3
       (.I0(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_5 ),
        .O(PSUM2__60_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_3__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_5 ),
        .O(PSUM2__60_carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_3__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_5 ),
        .O(PSUM2__60_carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_3__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_5 ),
        .O(PSUM2__60_carry_i_3__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_6 ),
        .O(PSUM2__60_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_6 ),
        .O(PSUM2__60_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_6 ),
        .O(PSUM2__60_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_6 ),
        .O(PSUM2__60_carry_i_4__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_5
       (.I0(\custom_alu/mult/mult16_3/PSUM2__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_7 ),
        .O(PSUM2__60_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_5__0
       (.I0(\custom_alu/mult/mult16_2/PSUM2__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_7 ),
        .O(PSUM2__60_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_5__1
       (.I0(\custom_alu/mult/mult16_1/PSUM2__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_7 ),
        .O(PSUM2__60_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM2__60_carry_i_5__2
       (.I0(\custom_alu/mult/mult16_0/PSUM2__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_7 ),
        .O(PSUM2__60_carry_i_5__2_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_1
       (.I0(ID_EX_Q[137]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[11]),
        .O(ALU_DIN1[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_10
       (.I0(ID_EX_Q[128]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[2]),
        .O(ALU_DIN1[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_11
       (.I0(ID_EX_Q[127]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[1]),
        .O(ALU_DIN1[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_12
       (.I0(ID_EX_Q[126]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[0]),
        .O(ALU_DIN1[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_2
       (.I0(ID_EX_Q[136]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[10]),
        .O(ALU_DIN1[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_3
       (.I0(ID_EX_Q[135]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[9]),
        .O(ALU_DIN1[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_4
       (.I0(ID_EX_Q[134]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[8]),
        .O(ALU_DIN1[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_5
       (.I0(ID_EX_Q[133]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[7]),
        .O(ALU_DIN1[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_6
       (.I0(ID_EX_Q[132]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[6]),
        .O(ALU_DIN1[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_7
       (.I0(ID_EX_Q[131]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[5]),
        .O(ALU_DIN1[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_8
       (.I0(ID_EX_Q[130]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[4]),
        .O(ALU_DIN1[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM2_i_9
       (.I0(ID_EX_Q[129]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[3]),
        .O(ALU_DIN1[3]));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_1
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[30]),
        .O(PSUM3__0_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_10
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM3__0_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_10__0
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM3__0_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_10__1
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM3__0_carry__0_i_10__1_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3__0_carry__0_i_10__2
       (.I0(ID_EX_Q[157]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[31]),
        .O(PSUM3__0_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_11
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM3__0_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_11__0
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[25]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[104]),
        .O(PSUM3__0_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_11__1
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM3__0_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_11__2
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[9]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[88]),
        .O(PSUM3__0_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_12
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM3__0_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_12__0
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[136]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM3__0_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_12__1
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM3__0_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__0_carry__0_i_12__2
       (.I0(ID_EX_Q[136]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[10]),
        .I3(ID_EX_Q[89]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[10]),
        .O(PSUM3__0_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__0_carry__0_i_13
       (.I0(ID_EX_Q[152]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[26]),
        .I3(ID_EX_Q[105]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[26]),
        .O(PSUM3__0_carry__0_i_13_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_1__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[14]),
        .O(PSUM3__0_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_1__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[30]),
        .O(PSUM3__0_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_1__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[14]),
        .O(PSUM3__0_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_2
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[29]),
        .O(PSUM3__0_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_2__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[13]),
        .O(PSUM3__0_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_2__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[29]),
        .O(PSUM3__0_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_2__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[13]),
        .O(PSUM3__0_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_3
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[28]),
        .O(PSUM3__0_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_3__0
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[12]),
        .O(PSUM3__0_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_3__1
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[12]),
        .O(PSUM3__0_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_3__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[28]),
        .O(PSUM3__0_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_4
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[27]),
        .O(PSUM3__0_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_4__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[11]),
        .O(PSUM3__0_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_4__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[27]),
        .O(PSUM3__0_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__0_i_4__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[11]),
        .O(PSUM3__0_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_5
       (.I0(PSUM3__0_carry__0_i_1_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM3__0_carry__0_i_9_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_5__0
       (.I0(PSUM3__0_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM3__0_carry__0_i_9__0_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_5__1
       (.I0(PSUM3__0_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM3__0_carry__0_i_9__1_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_5__2
       (.I0(PSUM3__0_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM3__0_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_6
       (.I0(PSUM3__0_carry__0_i_2_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM3__0_carry__0_i_11_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_6__0
       (.I0(PSUM3__0_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM3__0_carry__0_i_10_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_6__1
       (.I0(PSUM3__0_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM3__0_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_6__2
       (.I0(PSUM3__0_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM3__0_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_7
       (.I0(PSUM3__0_carry__0_i_3_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM3__0_carry__0_i_12_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM3__0_carry__0_i_7__0
       (.I0(PSUM3__0_carry__0_i_3__0_n_0),
        .I1(PSUM3__0_carry__0_i_11__2_n_0),
        .I2(ALU_DIN2[10]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM3__0_carry__0_i_7__1
       (.I0(PSUM3__0_carry__0_i_3__1_n_0),
        .I1(PSUM3__0_carry__0_i_11__0_n_0),
        .I2(ALU_DIN2[26]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_7__2
       (.I0(PSUM3__0_carry__0_i_3__2_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM3__0_carry__0_i_11__1_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_8
       (.I0(PSUM3__0_carry__0_i_4_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM3__0_carry__0_i_13_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_8__0
       (.I0(PSUM3__0_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM3__0_carry__0_i_12__2_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_8__1
       (.I0(PSUM3__0_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[25]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM3__0_carry__0_i_12__0_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__0_carry__0_i_8__2
       (.I0(PSUM3__0_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[9]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM3__0_carry__0_i_12__1_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_9
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM3__0_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_9__0
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[26]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[105]),
        .O(PSUM3__0_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_9__1
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM3__0_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry__0_i_9__2
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[10]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[89]),
        .O(PSUM3__0_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__0_carry__1_i_1
       (.I0(ID_EX_Q[105]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[26]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[25]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__0_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__0_carry__1_i_1__0
       (.I0(ID_EX_Q[105]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[26]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[25]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__0_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__0_carry__1_i_1__1
       (.I0(ID_EX_Q[89]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[10]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[9]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__0_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__0_carry__1_i_1__2
       (.I0(ID_EX_Q[89]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[10]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[9]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__0_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__1_i_2
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[24]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__0_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__1_i_2__0
       (.I0(ALU_DIN2[26]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[25]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__0_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__1_i_2__1
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[8]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__0_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__0_carry__1_i_2__2
       (.I0(ALU_DIN2[10]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[9]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__0_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__0_carry__1_i_3
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[26]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__0_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__0_carry__1_i_3__0
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__0_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__0_carry__1_i_3__1
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[88]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[10]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__0_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__0_carry__1_i_3__2
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[88]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[10]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__0_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__0_carry__1_i_4
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[26]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[25]),
        .O(PSUM3__0_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__0_carry__1_i_4__0
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[26]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[25]),
        .O(PSUM3__0_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__0_carry__1_i_4__1
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[10]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[9]),
        .O(PSUM3__0_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__0_carry__1_i_4__2
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[10]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[9]),
        .O(PSUM3__0_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_1
       (.I0(ALU_DIN2[25]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[26]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_1__0
       (.I0(ALU_DIN2[25]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[26]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[24]),
        .O(PSUM3__0_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_1__1
       (.I0(ALU_DIN2[9]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[10]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_1__2
       (.I0(ALU_DIN2[9]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[10]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[8]),
        .O(PSUM3__0_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h1DFFE200E200E200)) 
    PSUM3__0_carry_i_2
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__0_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h1DFFE200E200E200)) 
    PSUM3__0_carry_i_2__0
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[88]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[10]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__0_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__0_carry_i_2__1
       (.I0(ID_EX_Q[104]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[25]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__0_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__0_carry_i_2__2
       (.I0(ID_EX_Q[88]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[9]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[10]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__0_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__0_carry_i_3
       (.I0(ID_EX_Q[103]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[24]),
        .I3(ID_EX_Q[151]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[25]),
        .O(PSUM3__0_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__0_carry_i_3__0
       (.I0(ID_EX_Q[103]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[24]),
        .I3(ID_EX_Q[135]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[9]),
        .O(PSUM3__0_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__0_carry_i_3__1
       (.I0(ID_EX_Q[87]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[8]),
        .I3(ID_EX_Q[151]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[25]),
        .O(PSUM3__0_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__0_carry_i_3__2
       (.I0(ID_EX_Q[87]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[8]),
        .I3(ID_EX_Q[135]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[9]),
        .O(PSUM3__0_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__0_carry_i_4
       (.I0(ALU_DIN1[26]),
        .I1(PSUM3__0_carry_i_8_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[26]),
        .O(PSUM3__0_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__0_carry_i_4__0
       (.I0(ALU_DIN1[10]),
        .I1(PSUM3__0_carry_i_8__2_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[10]),
        .O(PSUM3__0_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__0_carry_i_4__1
       (.I0(ALU_DIN1[10]),
        .I1(PSUM3__0_carry_i_8__0_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[26]),
        .O(PSUM3__0_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__0_carry_i_4__2
       (.I0(ALU_DIN1[26]),
        .I1(PSUM3__0_carry_i_8__1_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[10]),
        .O(PSUM3__0_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_5
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[26]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[26]),
        .O(PSUM3__0_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_5__0
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[10]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[10]),
        .O(PSUM3__0_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_5__1
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[26]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[25]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[10]),
        .O(PSUM3__0_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__0_carry_i_5__2
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[10]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[9]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[26]),
        .O(PSUM3__0_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM3__0_carry_i_6
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[25]),
        .I2(ID_EX_Q[104]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[25]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__0_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM3__0_carry_i_6__0
       (.I0(ALU_DIN2[24]),
        .I1(ALU_DIN1[9]),
        .I2(ID_EX_Q[104]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[25]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__0_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM3__0_carry_i_6__1
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[25]),
        .I2(ID_EX_Q[88]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[9]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__0_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h7877788888888888)) 
    PSUM3__0_carry_i_6__2
       (.I0(ALU_DIN2[8]),
        .I1(ALU_DIN1[9]),
        .I2(ID_EX_Q[88]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[9]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__0_carry_i_6__2_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__0_carry_i_7
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM3__0_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__0_carry_i_7__0
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM3__0_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__0_carry_i_7__1
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM3__0_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__0_carry_i_7__2
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM3__0_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry_i_8
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM3__0_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry_i_8__0
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(EX_RF_RD2[24]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[103]),
        .O(PSUM3__0_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry_i_8__1
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM3__0_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__0_carry_i_8__2
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(EX_RF_RD2[8]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[87]),
        .O(PSUM3__0_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_1
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[30]),
        .O(PSUM3__30_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_10
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM3__30_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_10__0
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM3__30_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_10__1
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[154]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM3__30_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_10__2
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM3__30_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_11
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM3__30_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_11__0
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[138]),
        .I3(EX_RF_RD2[28]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[107]),
        .O(PSUM3__30_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_11__1
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM3__30_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__30_carry__0_i_11__2
       (.I0(ID_EX_Q[138]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[12]),
        .I3(ID_EX_Q[91]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[12]),
        .O(PSUM3__30_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_12
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM3__30_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_12__0
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[136]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM3__30_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_12__1
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM3__30_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_12__2
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[136]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM3__30_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_1__0
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[14]),
        .O(PSUM3__30_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_1__1
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[28]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[29]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[30]),
        .O(PSUM3__30_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_1__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[12]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[13]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[14]),
        .O(PSUM3__30_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_2
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[29]),
        .O(PSUM3__30_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_2__0
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[13]),
        .O(PSUM3__30_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_2__1
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[11]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[13]),
        .O(PSUM3__30_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_2__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[27]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[29]),
        .O(PSUM3__30_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_3
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[28]),
        .O(PSUM3__30_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_3__0
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[12]),
        .O(PSUM3__30_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_3__1
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[27]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[28]),
        .O(PSUM3__30_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_3__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[12]),
        .O(PSUM3__30_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_4
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[27]),
        .O(PSUM3__30_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_4__0
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[11]),
        .O(PSUM3__30_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_4__1
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[11]),
        .O(PSUM3__30_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__0_i_4__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[27]),
        .O(PSUM3__30_carry__0_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_5
       (.I0(PSUM3__30_carry__0_i_1_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM3__30_carry__0_i_9__1_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_5__0
       (.I0(PSUM3__30_carry__0_i_1__2_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM3__30_carry__0_i_9__2_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_5__1
       (.I0(PSUM3__30_carry__0_i_1__0_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[14]),
        .I3(PSUM3__30_carry__0_i_9_n_0),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_5__2
       (.I0(PSUM3__30_carry__0_i_1__1_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[30]),
        .I3(PSUM3__30_carry__0_i_9__0_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_6
       (.I0(PSUM3__30_carry__0_i_2_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM3__30_carry__0_i_10_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_6__0
       (.I0(PSUM3__30_carry__0_i_2__0_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM3__30_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_6__1
       (.I0(PSUM3__30_carry__0_i_2__1_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM3__30_carry__0_i_10__0_n_0),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_6__2
       (.I0(PSUM3__30_carry__0_i_2__2_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[29]),
        .I3(PSUM3__30_carry__0_i_10__1_n_0),
        .I4(ALU_DIN1[30]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_7
       (.I0(PSUM3__30_carry__0_i_3_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM3__30_carry__0_i_11_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM3__30_carry__0_i_7__0
       (.I0(PSUM3__30_carry__0_i_3__2_n_0),
        .I1(PSUM3__30_carry__0_i_11__2_n_0),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h9666699969996999)) 
    PSUM3__30_carry__0_i_7__1
       (.I0(PSUM3__30_carry__0_i_3__0_n_0),
        .I1(PSUM3__30_carry__0_i_11__0_n_0),
        .I2(ALU_DIN2[29]),
        .I3(ALU_DIN1[11]),
        .I4(ALU_DIN1[13]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_7__2
       (.I0(PSUM3__30_carry__0_i_3__1_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[28]),
        .I3(PSUM3__30_carry__0_i_11__1_n_0),
        .I4(ALU_DIN1[29]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_8
       (.I0(PSUM3__30_carry__0_i_4_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM3__30_carry__0_i_12_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_8__0
       (.I0(PSUM3__30_carry__0_i_4__0_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM3__30_carry__0_i_12__2_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_8__1
       (.I0(PSUM3__30_carry__0_i_4__1_n_0),
        .I1(ALU_DIN2[28]),
        .I2(ALU_DIN1[11]),
        .I3(PSUM3__30_carry__0_i_12__0_n_0),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry__0_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h956A6A956A956A95)) 
    PSUM3__30_carry__0_i_8__2
       (.I0(PSUM3__30_carry__0_i_4__2_n_0),
        .I1(ALU_DIN2[12]),
        .I2(ALU_DIN1[27]),
        .I3(PSUM3__30_carry__0_i_12__1_n_0),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_9
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[29]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[108]),
        .O(PSUM3__30_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry__0_i_9__0
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[13]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[92]),
        .O(PSUM3__30_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__30_carry__0_i_9__1
       (.I0(ID_EX_Q[155]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[29]),
        .I3(ID_EX_Q[108]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[29]),
        .O(PSUM3__30_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__30_carry__0_i_9__2
       (.I0(ID_EX_Q[139]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[13]),
        .I3(ID_EX_Q[92]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[13]),
        .O(PSUM3__30_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__30_carry__1_i_1
       (.I0(ID_EX_Q[108]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[29]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[28]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__30_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__30_carry__1_i_1__0
       (.I0(ID_EX_Q[108]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[29]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__30_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__30_carry__1_i_1__1
       (.I0(ID_EX_Q[92]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[13]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[12]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__30_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    PSUM3__30_carry__1_i_1__2
       (.I0(ID_EX_Q[92]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[13]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[12]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__30_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__1_i_2
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[27]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__30_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__1_i_2__0
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__30_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__1_i_2__1
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN2[28]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__30_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'hF888800080008000)) 
    PSUM3__30_carry__1_i_2__2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN2[12]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[11]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__30_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__30_carry__1_i_3
       (.I0(EX_RF_RD2[28]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[107]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[29]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__30_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__30_carry__1_i_3__0
       (.I0(EX_RF_RD2[28]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(ID_EX_Q[107]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[29]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__30_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__30_carry__1_i_3__1
       (.I0(EX_RF_RD2[12]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[91]),
        .I3(ALU_DIN1[30]),
        .I4(ALU_DIN2[13]),
        .I5(PSUM3__0_carry__0_i_10__2_n_0),
        .O(PSUM3__30_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h1DFF000000000000)) 
    PSUM3__30_carry__1_i_3__2
       (.I0(EX_RF_RD2[12]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[91]),
        .I3(ALU_DIN1[14]),
        .I4(ALU_DIN2[13]),
        .I5(ALU_DIN1[15]),
        .O(PSUM3__30_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__30_carry__1_i_4
       (.I0(ALU_DIN2[27]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[29]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[28]),
        .O(PSUM3__30_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__30_carry__1_i_4__0
       (.I0(ALU_DIN2[11]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[13]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[12]),
        .O(PSUM3__30_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__30_carry__1_i_4__1
       (.I0(ALU_DIN2[27]),
        .I1(ALU_DIN1[13]),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[29]),
        .I4(ALU_DIN1[15]),
        .I5(ALU_DIN2[28]),
        .O(PSUM3__30_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hE75F30007800F000)) 
    PSUM3__30_carry__1_i_4__2
       (.I0(ALU_DIN2[11]),
        .I1(ALU_DIN1[29]),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[13]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN2[12]),
        .O(PSUM3__30_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_1
       (.I0(ALU_DIN2[28]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[29]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_1__0
       (.I0(ALU_DIN2[12]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_1__1
       (.I0(ALU_DIN2[28]),
        .I1(ALU_DIN1[10]),
        .I2(ALU_DIN2[29]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN1[11]),
        .I5(ALU_DIN2[27]),
        .O(PSUM3__30_carry_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_1__2
       (.I0(ALU_DIN2[12]),
        .I1(ALU_DIN1[26]),
        .I2(ALU_DIN2[13]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN1[27]),
        .I5(ALU_DIN2[11]),
        .O(PSUM3__30_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_2
       (.I0(ID_EX_Q[107]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[28]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[29]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__30_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_2__0
       (.I0(ID_EX_Q[107]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[28]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[29]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__30_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_2__1
       (.I0(ID_EX_Q[91]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[12]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[13]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__30_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_2__2
       (.I0(ID_EX_Q[91]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[12]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[13]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__30_carry_i_2__2_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__30_carry_i_3
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ID_EX_Q[151]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[25]),
        .O(PSUM3__30_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__30_carry_i_3__0
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ID_EX_Q[135]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[9]),
        .O(PSUM3__30_carry_i_3__0_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__30_carry_i_3__1
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ID_EX_Q[151]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[25]),
        .O(PSUM3__30_carry_i_3__1_n_0));
  LUT6 #(
    .INIT(64'hB800B8B8B8000000)) 
    PSUM3__30_carry_i_3__2
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ID_EX_Q[135]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(EX_RF_RD1[9]),
        .O(PSUM3__30_carry_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__30_carry_i_4
       (.I0(ALU_DIN1[26]),
        .I1(PSUM3__30_carry_i_8__1_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[29]),
        .O(PSUM3__30_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__30_carry_i_4__0
       (.I0(ALU_DIN1[10]),
        .I1(PSUM3__30_carry_i_8__2_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[13]),
        .O(PSUM3__30_carry_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__30_carry_i_4__1
       (.I0(ALU_DIN1[10]),
        .I1(PSUM3__30_carry_i_8_n_0),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[29]),
        .O(PSUM3__30_carry_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h99C369C399339933)) 
    PSUM3__30_carry_i_4__2
       (.I0(ALU_DIN1[26]),
        .I1(PSUM3__30_carry_i_8__0_n_0),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[13]),
        .O(PSUM3__30_carry_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_5
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[29]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[26]),
        .O(PSUM3__30_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_5__0
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[29]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[28]),
        .I4(ALU_DIN2[27]),
        .I5(ALU_DIN1[10]),
        .O(PSUM3__30_carry_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_5__1
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN2[13]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[26]),
        .O(PSUM3__30_carry_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h8777788878887888)) 
    PSUM3__30_carry_i_5__2
       (.I0(ALU_DIN1[8]),
        .I1(ALU_DIN2[13]),
        .I2(ALU_DIN1[9]),
        .I3(ALU_DIN2[12]),
        .I4(ALU_DIN2[11]),
        .I5(ALU_DIN1[10]),
        .O(PSUM3__30_carry_i_5__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_6
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__30_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_6__0
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[28]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__30_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_6__1
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[12]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__30_carry_i_6__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B800B800)) 
    PSUM3__30_carry_i_6__2
       (.I0(ID_EX_Q[90]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[11]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[12]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__30_carry_i_6__2_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__30_carry_i_7
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM3__30_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__30_carry_i_7__0
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM3__30_carry_i_7__0_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__30_carry_i_7__1
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM3__30_carry_i_7__1_n_0));
  LUT6 #(
    .INIT(64'hE2E2E2000000E200)) 
    PSUM3__30_carry_i_7__2
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM3__30_carry_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry_i_8
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(EX_RF_RD2[27]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[106]),
        .O(PSUM3__30_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__30_carry_i_8__0
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[153]),
        .I3(EX_RF_RD2[11]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[90]),
        .O(PSUM3__30_carry_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__30_carry_i_8__1
       (.I0(ID_EX_Q[153]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[27]),
        .I3(ID_EX_Q[106]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[27]),
        .O(PSUM3__30_carry_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__30_carry_i_8__2
       (.I0(ID_EX_Q[137]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[11]),
        .I3(ID_EX_Q[90]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[11]),
        .O(PSUM3__30_carry_i_8__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__0_i_1
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM3__60_carry__0_i_9_n_0),
        .I5(PSUM3__60_carry__0_i_10_n_0),
        .O(PSUM3__60_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_10
       (.I0(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_7 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[25]),
        .O(PSUM3__60_carry__0_i_10_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_10__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_7 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[9]),
        .O(PSUM3__60_carry__0_i_10__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_10__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_7 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[25]),
        .O(PSUM3__60_carry__0_i_10__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_10__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_7 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[9]),
        .O(PSUM3__60_carry__0_i_10__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_11
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_7 ),
        .O(PSUM3__60_carry__0_i_11_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_11__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_7 ),
        .O(PSUM3__60_carry__0_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_11__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_7 ),
        .O(PSUM3__60_carry__0_i_11__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_11__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_6 ),
        .I5(\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_7 ),
        .O(PSUM3__60_carry__0_i_11__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_12
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[27]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_1 ),
        .O(PSUM3__60_carry__0_i_12_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_12__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[11]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_1 ),
        .O(PSUM3__60_carry__0_i_12__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_12__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[27]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_1 ),
        .O(PSUM3__60_carry__0_i_12__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_12__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[11]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_1 ),
        .O(PSUM3__60_carry__0_i_12__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_13
       (.I0(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_6 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[26]),
        .O(PSUM3__60_carry__0_i_13_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_13__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_6 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[10]),
        .O(PSUM3__60_carry__0_i_13__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_13__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_6 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[26]),
        .O(PSUM3__60_carry__0_i_13__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__0_i_13__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_6 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[10]),
        .O(PSUM3__60_carry__0_i_13__2_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM3__60_carry__0_i_14
       (.I0(ALU_DIN1[25]),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[30]),
        .I5(PSUM3__60_carry__0_i_11_n_0),
        .O(PSUM3__60_carry__0_i_14_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM3__60_carry__0_i_14__0
       (.I0(ALU_DIN1[9]),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[30]),
        .I5(PSUM3__60_carry__0_i_11__0_n_0),
        .O(PSUM3__60_carry__0_i_14__0_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM3__60_carry__0_i_14__1
       (.I0(ALU_DIN1[25]),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ),
        .I3(ALU_DIN1[26]),
        .I4(ALU_DIN2[14]),
        .I5(PSUM3__60_carry__0_i_11__1_n_0),
        .O(PSUM3__60_carry__0_i_14__1_n_0));
  LUT6 #(
    .INIT(64'h807FFFFF7F800000)) 
    PSUM3__60_carry__0_i_14__2
       (.I0(ALU_DIN1[9]),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ),
        .I2(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ),
        .I3(ALU_DIN1[10]),
        .I4(ALU_DIN2[14]),
        .I5(PSUM3__60_carry__0_i_11__2_n_0),
        .O(PSUM3__60_carry__0_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_15
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[24]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_4 ),
        .O(PSUM3__60_carry__0_i_15_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_15__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[8]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_4 ),
        .O(PSUM3__60_carry__0_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_15__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[24]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_4 ),
        .O(PSUM3__60_carry__0_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_15__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[8]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_7 ),
        .I5(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_4 ),
        .O(PSUM3__60_carry__0_i_15__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__0_i_1__0
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM3__60_carry__0_i_9__0_n_0),
        .I5(PSUM3__60_carry__0_i_10__0_n_0),
        .O(PSUM3__60_carry__0_i_1__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__0_i_1__1
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM3__60_carry__0_i_9__1_n_0),
        .I5(PSUM3__60_carry__0_i_10__1_n_0),
        .O(PSUM3__60_carry__0_i_1__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__0_i_1__2
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM3__60_carry__0_i_9__2_n_0),
        .I5(PSUM3__60_carry__0_i_10__2_n_0),
        .O(PSUM3__60_carry__0_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM3__60_carry__0_i_2
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[26]),
        .I2(PSUM3__60_carry__0_i_11_n_0),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM3__60_carry__0_i_2__0
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[10]),
        .I2(PSUM3__60_carry__0_i_11__0_n_0),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM3__60_carry__0_i_2__1
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[26]),
        .I2(PSUM3__60_carry__0_i_11__1_n_0),
        .I3(ALU_DIN1[25]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h8A08080808080808)) 
    PSUM3__60_carry__0_i_2__2
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[10]),
        .I2(PSUM3__60_carry__0_i_11__2_n_0),
        .I3(ALU_DIN1[9]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ),
        .I5(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM3__60_carry__0_i_3
       (.I0(PSUM3__60_carry__0_i_11_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN1[26]),
        .I3(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ),
        .I5(ALU_DIN1[25]),
        .O(PSUM3__60_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM3__60_carry__0_i_3__0
       (.I0(PSUM3__60_carry__0_i_11__0_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN1[10]),
        .I3(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ),
        .I5(ALU_DIN1[9]),
        .O(PSUM3__60_carry__0_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM3__60_carry__0_i_3__1
       (.I0(PSUM3__60_carry__0_i_11__1_n_0),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN1[26]),
        .I3(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ),
        .I5(ALU_DIN1[25]),
        .O(PSUM3__60_carry__0_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h5995959595959595)) 
    PSUM3__60_carry__0_i_3__2
       (.I0(PSUM3__60_carry__0_i_11__2_n_0),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN1[10]),
        .I3(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ),
        .I5(ALU_DIN1[9]),
        .O(PSUM3__60_carry__0_i_3__2_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM3__60_carry__0_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_7 ),
        .I2(ALU_DIN1[24]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM3__60_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM3__60_carry__0_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_7 ),
        .I2(ALU_DIN1[8]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM3__60_carry__0_i_4__0_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM3__60_carry__0_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_7 ),
        .I2(ALU_DIN1[24]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM3__60_carry__0_i_4__1_n_0));
  LUT6 #(
    .INIT(64'h9696966666669666)) 
    PSUM3__60_carry__0_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_7 ),
        .I2(ALU_DIN1[8]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM3__60_carry__0_i_4__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_5
       (.I0(PSUM3__60_carry__0_i_1_n_0),
        .I1(PSUM3__60_carry__0_i_12_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM3__60_carry__0_i_13_n_0),
        .O(PSUM3__60_carry__0_i_5_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_5__0
       (.I0(PSUM3__60_carry__0_i_1__0_n_0),
        .I1(PSUM3__60_carry__0_i_12__0_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM3__60_carry__0_i_13__0_n_0),
        .O(PSUM3__60_carry__0_i_5__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_5__1
       (.I0(PSUM3__60_carry__0_i_1__1_n_0),
        .I1(PSUM3__60_carry__0_i_12__1_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM3__60_carry__0_i_13__1_n_0),
        .O(PSUM3__60_carry__0_i_5__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_5__2
       (.I0(PSUM3__60_carry__0_i_1__2_n_0),
        .I1(PSUM3__60_carry__0_i_12__2_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM3__60_carry__0_i_13__2_n_0),
        .O(PSUM3__60_carry__0_i_5__2_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_6
       (.I0(PSUM3__60_carry__0_i_2_n_0),
        .I1(PSUM3__60_carry__0_i_9_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM3__60_carry__0_i_10_n_0),
        .O(PSUM3__60_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_6__0
       (.I0(PSUM3__60_carry__0_i_2__0_n_0),
        .I1(PSUM3__60_carry__0_i_9__0_n_0),
        .I2(ALU_DIN2[30]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM3__60_carry__0_i_10__0_n_0),
        .O(PSUM3__60_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_6__1
       (.I0(PSUM3__60_carry__0_i_2__1_n_0),
        .I1(PSUM3__60_carry__0_i_9__1_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM3__60_carry__0_i_10__1_n_0),
        .O(PSUM3__60_carry__0_i_6__1_n_0));
  LUT5 #(
    .INIT(32'h96666999)) 
    PSUM3__60_carry__0_i_6__2
       (.I0(PSUM3__60_carry__0_i_2__2_n_0),
        .I1(PSUM3__60_carry__0_i_9__2_n_0),
        .I2(ALU_DIN2[14]),
        .I3(ALU_DIN1[11]),
        .I4(PSUM3__60_carry__0_i_10__2_n_0),
        .O(PSUM3__60_carry__0_i_6__2_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM3__60_carry__0_i_7
       (.I0(PSUM3__60_carry__0_i_14_n_0),
        .I1(ALU_DIN1[24]),
        .I2(ALU_DIN2[31]),
        .I3(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_7 ),
        .O(PSUM3__60_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM3__60_carry__0_i_7__0
       (.I0(PSUM3__60_carry__0_i_14__0_n_0),
        .I1(ALU_DIN1[8]),
        .I2(ALU_DIN2[31]),
        .I3(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_7 ),
        .O(PSUM3__60_carry__0_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM3__60_carry__0_i_7__1
       (.I0(PSUM3__60_carry__0_i_14__1_n_0),
        .I1(ALU_DIN1[24]),
        .I2(ALU_DIN2[15]),
        .I3(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_7 ),
        .O(PSUM3__60_carry__0_i_7__1_n_0));
  LUT5 #(
    .INIT(32'hAA959555)) 
    PSUM3__60_carry__0_i_7__2
       (.I0(PSUM3__60_carry__0_i_14__2_n_0),
        .I1(ALU_DIN1[8]),
        .I2(ALU_DIN2[15]),
        .I3(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_7 ),
        .O(PSUM3__60_carry__0_i_7__2_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM3__60_carry__0_i_8
       (.I0(PSUM3__60_carry__0_i_15_n_0),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[30]),
        .I3(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_8_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM3__60_carry__0_i_8__0
       (.I0(PSUM3__60_carry__0_i_15__0_n_0),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[30]),
        .I3(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM3__60_carry__0_i_8__1
       (.I0(PSUM3__60_carry__0_i_15__1_n_0),
        .I1(ALU_DIN1[25]),
        .I2(ALU_DIN2[14]),
        .I3(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_8__1_n_0));
  LUT5 #(
    .INIT(32'h6A959595)) 
    PSUM3__60_carry__0_i_8__2
       (.I0(PSUM3__60_carry__0_i_15__2_n_0),
        .I1(ALU_DIN1[9]),
        .I2(ALU_DIN2[14]),
        .I3(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ),
        .I4(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ),
        .O(PSUM3__60_carry__0_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_9
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[26]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_6 ),
        .O(PSUM3__60_carry__0_i_9_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_9__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[10]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_6 ),
        .O(PSUM3__60_carry__0_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_9__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[26]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_6 ),
        .O(PSUM3__60_carry__0_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h47FFB800B80047FF)) 
    PSUM3__60_carry__0_i_9__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[10]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_5 ),
        .I5(\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_6 ),
        .O(PSUM3__60_carry__0_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_1
       (.I0(PSUM3__60_carry__1_i_9_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_6 ),
        .I5(ALU_DIN1[29]),
        .O(PSUM3__60_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_10
       (.I0(EX_RF_RD1[14]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[140]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM3__60_carry__1_i_10_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_10__0
       (.I0(EX_RF_RD1[30]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[156]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM3__60_carry__1_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__60_carry__1_i_10__1
       (.I0(ID_EX_Q[156]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[30]),
        .I3(ID_EX_Q[109]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[30]),
        .O(PSUM3__60_carry__1_i_10__1_n_0));
  LUT6 #(
    .INIT(64'h47FF474747FFFFFF)) 
    PSUM3__60_carry__1_i_10__2
       (.I0(ID_EX_Q[140]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(EX_RF_RD1[14]),
        .I3(ID_EX_Q[93]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[14]),
        .O(PSUM3__60_carry__1_i_10__2_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__1_i_11
       (.I0(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_1 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[27]),
        .O(PSUM3__60_carry__1_i_11_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__1_i_11__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_1 ),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I4(EX_RF_RD2[31]),
        .I5(ALU_DIN1[11]),
        .O(PSUM3__60_carry__1_i_11__0_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__1_i_11__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_1 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[27]),
        .O(PSUM3__60_carry__1_i_11__1_n_0));
  LUT6 #(
    .INIT(64'hE8EEE88888888888)) 
    PSUM3__60_carry__1_i_11__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_1 ),
        .I2(ID_EX_Q[94]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[15]),
        .I5(ALU_DIN1[11]),
        .O(PSUM3__60_carry__1_i_11__2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM3__60_carry__1_i_12
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM3__60_carry__1_i_12__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_12__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM3__60_carry__1_i_12__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_12__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'h47FFFFFF)) 
    PSUM3__60_carry__1_i_12__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_12__2_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_13
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[30]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_13__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[14]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_13__0_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_13__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[30]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_13__1_n_0));
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_13__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[14]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_13__2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_14
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_14_n_0));
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_14__0
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_14__0_n_0));
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_14__1
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[29]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_14__1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'hB80047FF)) 
    PSUM3__60_carry__1_i_14__2
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[15]),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_14__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_15
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM3__60_carry__1_i_15_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_15__0
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM3__60_carry__1_i_15__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_15__1
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[155]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM3__60_carry__1_i_15__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_15__2
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[139]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM3__60_carry__1_i_15__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_1__0
       (.I0(PSUM3__60_carry__1_i_9__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_6 ),
        .I5(ALU_DIN1[13]),
        .O(PSUM3__60_carry__1_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_1__1
       (.I0(PSUM3__60_carry__1_i_9__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_6 ),
        .I5(ALU_DIN1[29]),
        .O(PSUM3__60_carry__1_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_1__2
       (.I0(PSUM3__60_carry__1_i_9__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_6 ),
        .I5(ALU_DIN1[13]),
        .O(PSUM3__60_carry__1_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_2
       (.I0(PSUM3__60_carry__1_i_10__1_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_6 ),
        .I2(ALU_DIN1[29]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_7 ),
        .I5(ALU_DIN1[28]),
        .O(PSUM3__60_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_2__0
       (.I0(PSUM3__60_carry__1_i_10__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_6 ),
        .I2(ALU_DIN1[13]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_7 ),
        .I5(ALU_DIN1[12]),
        .O(PSUM3__60_carry__1_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_2__1
       (.I0(PSUM3__60_carry__1_i_10_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_6 ),
        .I2(ALU_DIN1[13]),
        .I3(ALU_DIN2[31]),
        .I4(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_7 ),
        .I5(ALU_DIN1[12]),
        .O(PSUM3__60_carry__1_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h7D44144414441444)) 
    PSUM3__60_carry__1_i_2__2
       (.I0(PSUM3__60_carry__1_i_10__0_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_6 ),
        .I2(ALU_DIN1[29]),
        .I3(ALU_DIN2[15]),
        .I4(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_7 ),
        .I5(ALU_DIN1[28]),
        .O(PSUM3__60_carry__1_i_2__2_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM3__60_carry__1_i_3
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[29]),
        .I2(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_7 ),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[31]),
        .I5(PSUM3__60_carry__1_i_11_n_0),
        .O(PSUM3__60_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM3__60_carry__1_i_3__0
       (.I0(ALU_DIN2[30]),
        .I1(ALU_DIN1[13]),
        .I2(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_7 ),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[31]),
        .I5(PSUM3__60_carry__1_i_11__0_n_0),
        .O(PSUM3__60_carry__1_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM3__60_carry__1_i_3__1
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[29]),
        .I2(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_7 ),
        .I3(ALU_DIN1[28]),
        .I4(ALU_DIN2[15]),
        .I5(PSUM3__60_carry__1_i_11__1_n_0),
        .O(PSUM3__60_carry__1_i_3__1_n_0));
  LUT6 #(
    .INIT(64'h8FF8F8F808808080)) 
    PSUM3__60_carry__1_i_3__2
       (.I0(ALU_DIN2[14]),
        .I1(ALU_DIN1[13]),
        .I2(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_7 ),
        .I3(ALU_DIN1[12]),
        .I4(ALU_DIN2[15]),
        .I5(PSUM3__60_carry__1_i_11__2_n_0),
        .O(PSUM3__60_carry__1_i_3__2_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__1_i_4
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM3__60_carry__0_i_12_n_0),
        .I5(PSUM3__60_carry__0_i_13_n_0),
        .O(PSUM3__60_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__1_i_4__0
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM3__60_carry__0_i_12__0_n_0),
        .I5(PSUM3__60_carry__0_i_13__0_n_0),
        .O(PSUM3__60_carry__1_i_4__0_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__1_i_4__1
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[28]),
        .I4(PSUM3__60_carry__0_i_12__1_n_0),
        .I5(PSUM3__60_carry__0_i_13__1_n_0),
        .O(PSUM3__60_carry__1_i_4__1_n_0));
  LUT6 #(
    .INIT(64'hB800FFFF0000B800)) 
    PSUM3__60_carry__1_i_4__2
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[14]),
        .I3(ALU_DIN1[12]),
        .I4(PSUM3__60_carry__0_i_12__2_n_0),
        .I5(PSUM3__60_carry__0_i_13__2_n_0),
        .O(PSUM3__60_carry__1_i_4__2_n_0));
  LUT6 #(
    .INIT(64'h4DF52D552450B400)) 
    PSUM3__60_carry__1_i_5
       (.I0(PSUM3__60_carry__1_i_12_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN2[31]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[30]),
        .I5(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_5_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM3__60_carry__1_i_5__0
       (.I0(PSUM3__60_carry__1_i_12__2_n_0),
        .I1(ALU_DIN2[14]),
        .I2(ALU_DIN1[15]),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[14]),
        .I5(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_5__0_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM3__60_carry__1_i_5__1
       (.I0(PSUM3__60_carry__1_i_12__0_n_0),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN1[15]),
        .I3(ALU_DIN2[31]),
        .I4(ALU_DIN1[14]),
        .I5(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_5__1_n_0));
  LUT6 #(
    .INIT(64'h4FD525D52540B040)) 
    PSUM3__60_carry__1_i_5__2
       (.I0(PSUM3__60_carry__1_i_12__1_n_0),
        .I1(ALU_DIN2[14]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[30]),
        .I5(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_1 ),
        .O(PSUM3__60_carry__1_i_5__2_n_0));
  LUT5 #(
    .INIT(32'h69999666)) 
    PSUM3__60_carry__1_i_6
       (.I0(PSUM3__60_carry__1_i_2_n_0),
        .I1(PSUM3__60_carry__1_i_13_n_0),
        .I2(ALU_DIN2[30]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(PSUM3__60_carry__1_i_12_n_0),
        .O(PSUM3__60_carry__1_i_6_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM3__60_carry__1_i_6__0
       (.I0(PSUM3__60_carry__1_i_2__0_n_0),
        .I1(PSUM3__60_carry__1_i_13__2_n_0),
        .I2(PSUM3__60_carry__1_i_9__2_n_0),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[13]),
        .I5(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM3__60_carry__1_i_6__1
       (.I0(PSUM3__60_carry__1_i_2__1_n_0),
        .I1(PSUM3__60_carry__1_i_13__0_n_0),
        .I2(PSUM3__60_carry__1_i_9__0_n_0),
        .I3(ALU_DIN2[31]),
        .I4(ALU_DIN1[13]),
        .I5(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_6 ),
        .O(PSUM3__60_carry__1_i_6__1_n_0));
  LUT5 #(
    .INIT(32'h69999666)) 
    PSUM3__60_carry__1_i_6__2
       (.I0(PSUM3__60_carry__1_i_2__2_n_0),
        .I1(PSUM3__60_carry__1_i_13__1_n_0),
        .I2(ALU_DIN2[14]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(PSUM3__60_carry__1_i_12__1_n_0),
        .O(PSUM3__60_carry__1_i_6__2_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM3__60_carry__1_i_7
       (.I0(PSUM3__60_carry__1_i_3_n_0),
        .I1(PSUM3__60_carry__1_i_14_n_0),
        .I2(PSUM3__60_carry__1_i_10__1_n_0),
        .I3(ALU_DIN2[31]),
        .I4(ALU_DIN1[28]),
        .I5(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_7 ),
        .O(PSUM3__60_carry__1_i_7_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM3__60_carry__1_i_7__0
       (.I0(PSUM3__60_carry__1_i_3__2_n_0),
        .I1(PSUM3__60_carry__1_i_14__2_n_0),
        .I2(PSUM3__60_carry__1_i_10__2_n_0),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[12]),
        .I5(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_7 ),
        .O(PSUM3__60_carry__1_i_7__0_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM3__60_carry__1_i_7__1
       (.I0(PSUM3__60_carry__1_i_3__0_n_0),
        .I1(PSUM3__60_carry__1_i_14__0_n_0),
        .I2(PSUM3__60_carry__1_i_10_n_0),
        .I3(ALU_DIN2[31]),
        .I4(ALU_DIN1[12]),
        .I5(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_7 ),
        .O(PSUM3__60_carry__1_i_7__1_n_0));
  LUT6 #(
    .INIT(64'h6996969696969696)) 
    PSUM3__60_carry__1_i_7__2
       (.I0(PSUM3__60_carry__1_i_3__1_n_0),
        .I1(PSUM3__60_carry__1_i_14__1_n_0),
        .I2(PSUM3__60_carry__1_i_10__0_n_0),
        .I3(ALU_DIN2[15]),
        .I4(ALU_DIN1[28]),
        .I5(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_7 ),
        .O(PSUM3__60_carry__1_i_7__2_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM3__60_carry__1_i_8
       (.I0(PSUM3__60_carry__1_i_4_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_7 ),
        .I2(ALU_DIN1[28]),
        .I3(ALU_DIN2[31]),
        .I4(PSUM3__60_carry__1_i_15_n_0),
        .I5(PSUM3__60_carry__1_i_11_n_0),
        .O(PSUM3__60_carry__1_i_8_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM3__60_carry__1_i_8__0
       (.I0(PSUM3__60_carry__1_i_4__0_n_0),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_7 ),
        .I2(ALU_DIN1[12]),
        .I3(ALU_DIN2[31]),
        .I4(PSUM3__60_carry__1_i_15__0_n_0),
        .I5(PSUM3__60_carry__1_i_11__0_n_0),
        .O(PSUM3__60_carry__1_i_8__0_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM3__60_carry__1_i_8__1
       (.I0(PSUM3__60_carry__1_i_4__1_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_7 ),
        .I2(ALU_DIN1[28]),
        .I3(ALU_DIN2[15]),
        .I4(PSUM3__60_carry__1_i_15__1_n_0),
        .I5(PSUM3__60_carry__1_i_11__1_n_0),
        .O(PSUM3__60_carry__1_i_8__1_n_0));
  LUT6 #(
    .INIT(64'h6999966696666999)) 
    PSUM3__60_carry__1_i_8__2
       (.I0(PSUM3__60_carry__1_i_4__2_n_0),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_7 ),
        .I2(ALU_DIN1[12]),
        .I3(ALU_DIN2[15]),
        .I4(PSUM3__60_carry__1_i_15__2_n_0),
        .I5(PSUM3__60_carry__1_i_11__2_n_0),
        .O(PSUM3__60_carry__1_i_8__2_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_9
       (.I0(EX_RF_RD1[31]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[157]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM3__60_carry__1_i_9_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_9__0
       (.I0(EX_RF_RD1[15]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I2(ID_EX_Q[141]),
        .I3(EX_RF_RD2[30]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__0_n_0 ),
        .I5(ID_EX_Q[109]),
        .O(PSUM3__60_carry__1_i_9__0_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_9__1
       (.I0(EX_RF_RD1[31]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[157]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__1_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM3__60_carry__1_i_9__1_n_0));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF)) 
    PSUM3__60_carry__1_i_9__2
       (.I0(EX_RF_RD1[15]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I2(ID_EX_Q[141]),
        .I3(EX_RF_RD2[14]),
        .I4(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I5(ID_EX_Q[93]),
        .O(PSUM3__60_carry__1_i_9__2_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM3__60_carry__2_i_1
       (.I0(PSUM3__0_carry__0_i_10__2_n_0),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM3__60_carry__2_i_1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM3__60_carry__2_i_1__0
       (.I0(ALU_DIN1[15]),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM3__60_carry__2_i_1__0_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM3__60_carry__2_i_1__1
       (.I0(ALU_DIN1[15]),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[14]),
        .I3(EX_RF_RD2[31]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[110]),
        .O(PSUM3__60_carry__2_i_1__1_n_0));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    PSUM3__60_carry__2_i_1__2
       (.I0(PSUM3__0_carry__0_i_10__2_n_0),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_1 ),
        .I2(ALU_DIN1[30]),
        .I3(EX_RF_RD2[15]),
        .I4(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I5(ID_EX_Q[94]),
        .O(PSUM3__60_carry__2_i_1__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_1
       (.I0(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ),
        .O(PSUM3__60_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_1__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ),
        .O(PSUM3__60_carry_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_1__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ),
        .O(PSUM3__60_carry_i_1__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_1__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ),
        .O(PSUM3__60_carry_i_1__2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM3__60_carry_i_2
       (.I0(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ),
        .I2(ID_EX_Q[109]),
        .I3(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I4(EX_RF_RD2[30]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__60_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM3__60_carry_i_2__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ),
        .I2(ID_EX_Q[109]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[30]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__60_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM3__60_carry_i_2__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ),
        .I2(ID_EX_Q[93]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[14]),
        .I5(ALU_DIN1[24]),
        .O(PSUM3__60_carry_i_2__1_n_0));
  LUT6 #(
    .INIT(64'h9699966666666666)) 
    PSUM3__60_carry_i_2__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ),
        .I2(ID_EX_Q[93]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[14]),
        .I5(ALU_DIN1[8]),
        .O(PSUM3__60_carry_i_2__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_3
       (.I0(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_5 ),
        .O(PSUM3__60_carry_i_3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_3__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_5 ),
        .O(PSUM3__60_carry_i_3__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_3__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_5 ),
        .O(PSUM3__60_carry_i_3__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_3__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_6 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_5 ),
        .O(PSUM3__60_carry_i_3__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_4
       (.I0(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_6 ),
        .O(PSUM3__60_carry_i_4_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_4__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_6 ),
        .O(PSUM3__60_carry_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_4__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_6 ),
        .O(PSUM3__60_carry_i_4__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_4__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_7 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_6 ),
        .O(PSUM3__60_carry_i_4__2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_5
       (.I0(\custom_alu/mult/mult16_3/PSUM3__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_7 ),
        .O(PSUM3__60_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_5__0
       (.I0(\custom_alu/mult/mult16_2/PSUM3__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_7 ),
        .O(PSUM3__60_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_5__1
       (.I0(\custom_alu/mult/mult16_1/PSUM3__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_7 ),
        .O(PSUM3__60_carry_i_5__1_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    PSUM3__60_carry_i_5__2
       (.I0(\custom_alu/mult/mult16_0/PSUM3__0_carry_n_4 ),
        .I1(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_7 ),
        .O(PSUM3__60_carry_i_5__2_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    PSUM3_i_1
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN2[30]),
        .I2(ALU_DIN2[27]),
        .I3(ALU_DIN2[28]),
        .I4(PSUM3_i_25_n_0),
        .O(\custom_alu/fp32_mult/op_b1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_10
       (.I0(ID_EX_Q[93]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[14]),
        .O(ALU_DIN2[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_11
       (.I0(ID_EX_Q[92]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[13]),
        .O(ALU_DIN2[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_12
       (.I0(ID_EX_Q[91]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[12]),
        .O(ALU_DIN2[12]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    PSUM3_i_13
       (.I0(ALU_DIN1[26]),
        .I1(ALU_DIN1[30]),
        .I2(ALU_DIN1[25]),
        .I3(ALU_DIN1[27]),
        .I4(PSUM3_i_26_n_0),
        .O(\custom_alu/fp32_mult/op_a1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_14
       (.I0(ID_EX_Q[148]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[22]),
        .O(ALU_DIN1[22]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_15
       (.I0(ID_EX_Q[147]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[21]),
        .O(ALU_DIN1[21]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_16
       (.I0(ID_EX_Q[146]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[20]),
        .O(ALU_DIN1[20]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_17
       (.I0(ID_EX_Q[145]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[19]),
        .O(ALU_DIN1[19]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_18
       (.I0(ID_EX_Q[144]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[18]),
        .O(ALU_DIN1[18]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_19
       (.I0(ID_EX_Q[143]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[17]),
        .O(ALU_DIN1[17]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_2
       (.I0(ID_EX_Q[101]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[22]),
        .O(ALU_DIN2[22]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_20
       (.I0(ID_EX_Q[142]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[16]),
        .O(ALU_DIN1[16]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_21
       (.I0(ID_EX_Q[141]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[15]),
        .O(ALU_DIN1[15]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_22
       (.I0(ID_EX_Q[140]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[14]),
        .O(ALU_DIN1[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_23
       (.I0(ID_EX_Q[139]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[13]),
        .O(ALU_DIN1[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_24
       (.I0(ID_EX_Q[138]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[12]),
        .O(ALU_DIN1[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEA)) 
    PSUM3_i_25
       (.I0(ALU_DIN2[24]),
        .I1(ID_EX_Q[102]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[23]),
        .I4(ALU_DIN2[26]),
        .I5(ALU_DIN2[25]),
        .O(PSUM3_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFEFEFE)) 
    PSUM3_i_26
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN1[23]),
        .I2(ALU_DIN1[29]),
        .I3(ID_EX_Q[154]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I5(EX_RF_RD1[28]),
        .O(PSUM3_i_26_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_3
       (.I0(ID_EX_Q[100]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[21]),
        .O(ALU_DIN2[21]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_4
       (.I0(ID_EX_Q[99]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[20]),
        .O(ALU_DIN2[20]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_5
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[19]),
        .O(ALU_DIN2[19]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_6
       (.I0(ID_EX_Q[97]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[18]),
        .O(ALU_DIN2[18]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_7
       (.I0(ID_EX_Q[96]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[17]),
        .O(ALU_DIN2[17]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_8
       (.I0(ID_EX_Q[95]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[16]),
        .O(ALU_DIN2[16]));
  LUT3 #(
    .INIT(8'hB8)) 
    PSUM3_i_9
       (.I0(ID_EX_Q[94]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[15]),
        .O(ALU_DIN2[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAAAE)) 
    \Q[0]_i_1 
       (.I0(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .I1(\Q[0]_i_3_n_0 ),
        .I2(\Q[160]_i_2_n_0 ),
        .I3(I_MEM_DOUT_FILTERED[4]),
        .I4(CUSTOM_INSTRUCTION_STALL_CYCLE[2]),
        .I5(\Q[27]_i_2_n_0 ),
        .O(CUSTOM_EN));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0100)) 
    \Q[0]_i_1__0 
       (.I0(\Q[160]_i_2_n_0 ),
        .I1(I_MEM_DOUT_FILTERED[4]),
        .I2(I_MEM_DOUT_FILTERED[5]),
        .I3(\Q[0]_i_3_n_0 ),
        .I4(CUSTOM_ALU_SEL[26]),
        .I5(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .O(CUSTOM_RD));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \Q[0]_i_1__1 
       (.I0(I_MEM_DOUT_IBUF[3]),
        .I1(I_MEM_DOUT_IBUF[4]),
        .I2(I_MEM_DOUT_IBUF[5]),
        .I3(I_MEM_DOUT_IBUF[6]),
        .I4(EX_BR_TAKEN),
        .I5(I_MEM_DOUT_IBUF[2]),
        .O(DECODED_INSTRUCTION[12]));
  LUT6 #(
    .INIT(64'h00000000EE2E2222)) 
    \Q[0]_i_1__2 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[1] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/sel0 [23]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [0]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[0]_i_1__3 
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[31]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .O(\custom_alu/fp32_add/p_1_in ));
  LUT5 #(
    .INIT(32'hFFE400E4)) 
    \Q[0]_i_1__4 
       (.I0(EX_BR_TAKEN),
        .I1(\FF_IF_ID_PCADD/Q_reg_n_0_[0] ),
        .I2(IF_PC2[0]),
        .I3(STALL_EN),
        .I4(ID_PC[0]),
        .O(\Q[0]_i_1__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[0]_i_1__5 
       (.I0(I_MEM_DOUT_IBUF[7]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[7]));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \Q[0]_i_1__6 
       (.I0(STALL_COUNTER_D1),
        .I1(STALL_COUNTER_Q[0]),
        .O(STALL_COUNTER_D[0]));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \Q[0]_i_2 
       (.I0(I_MEM_DOUT_IBUF[14]),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(\Q[31]_i_2_n_0 ),
        .O(CUSTOM_INSTRUCTION_STALL_CYCLE[2]));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \Q[0]_i_2__0 
       (.I0(EX_BR_TAKEN),
        .I1(I_MEM_DOUT_IBUF[4]),
        .O(I_MEM_DOUT_FILTERED[4]));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \Q[0]_i_3 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[6]),
        .I2(EX_BR_TAKEN),
        .I3(I_MEM_DOUT_IBUF[3]),
        .O(\Q[0]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[100]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(CRF_RA2_OBUF[1]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[21]));
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[101]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(CRF_RA2_OBUF[2]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[22]));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[102]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(CRF_RA2_OBUF[3]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[23]));
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[103]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(CRF_RA2_OBUF[4]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[24]));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[104]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[25]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[25]));
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[105]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[26]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[26]));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[106]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[27]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[27]));
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[107]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[28]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[28]));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[108]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[29]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[29]));
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[109]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[30]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[30]));
  LUT6 #(
    .INIT(64'hAAAAAAAAEEE2FFFF)) 
    \Q[109]_i_2 
       (.I0(\Q[109]_i_3_n_0 ),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[4]),
        .I5(EX_BR_TAKEN),
        .O(\Q[109]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT4 #(
    .INIT(16'hFFFD)) 
    \Q[109]_i_3 
       (.I0(I_MEM_DOUT_IBUF[12]),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[5]),
        .I3(EX_BR_TAKEN),
        .O(\Q[109]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[10]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [10]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [9]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [10]));
  LUT5 #(
    .INIT(32'h0000EEF0)) 
    \Q[10]_i_1__0 
       (.I0(\Q[10]_i_2_n_0 ),
        .I1(\Q[10]_i_3__1_n_0 ),
        .I2(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[11] ),
        .I3(\Q[30]_i_2__1_n_0 ),
        .I4(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [10]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[10]_i_1__1 
       (.I0(\Q[10]_i_2__0_n_0 ),
        .I1(\Q[10]_i_3_n_0 ),
        .I2(\Q[10]_i_4_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[5]),
        .O(data0[5]));
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \Q[10]_i_1__2 
       (.I0(\Q[10]_i_2__1_n_0 ),
        .I1(\Q[11]_i_3__0_n_0 ),
        .I2(\Q[10]_i_3__0_n_0 ),
        .I3(\Q[11]_i_5__1_n_0 ),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(EX_MEM_Q[10]),
        .O(data1[5]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[10]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [10]),
        .O(\Q[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[10]_i_2__0 
       (.I0(\custom_alu/MULT [5]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [37]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [5]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[10]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[10]_i_2__1 
       (.I0(D_MEM_DOUT_IBUF[13]),
        .I1(D_MEM_DOUT_IBUF[5]),
        .I2(D_MEM_DOUT_IBUF[29]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[21]),
        .O(\Q[10]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \Q[10]_i_3 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [5]),
        .O(\Q[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[10]_i_3__0 
       (.I0(D_MEM_DOUT_IBUF[5]),
        .I1(D_MEM_DOUT_IBUF[21]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[29]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[13]),
        .O(\Q[10]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h00F80000)) 
    \Q[10]_i_3__1 
       (.I0(\custom_alu/fp32_add/sel0 [9]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\Q[10]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [23]),
        .I4(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[10]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000032330233)) 
    \Q[10]_i_4 
       (.I0(INT0_carry__0_i_9_n_0),
        .I1(EX_CUSTOM_ALU_SEL[28]),
        .I2(ALU_DIN1[31]),
        .I3(EX_CUSTOM_ALU_SEL[27]),
        .I4(\custom_alu/fp2int/INT0 [5]),
        .I5(\Q[52]_i_5_n_0 ),
        .O(\Q[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5555510100005101)) 
    \Q[10]_i_4__0 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .I1(\Q[10]_i_5_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [7]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [8]),
        .O(\Q[10]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[10]_i_5 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [5]),
        .I3(\custom_alu/fp32_add/sel0 [18]),
        .I4(\Q[10]_i_6_n_0 ),
        .O(\Q[10]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h5555303F)) 
    \Q[10]_i_6 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [3]),
        .I2(\custom_alu/fp32_add/sel0 [16]),
        .I3(\Q[10]_i_7_n_0 ),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[10]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [13]),
        .O(\Q[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCCCCCCCCCCC8C)) 
    \Q[110]_i_1 
       (.I0(\Q[123]_i_3_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[12]),
        .I3(I_MEM_DOUT_IBUF[13]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(EX_BR_TAKEN),
        .O(ID_IMMEDIATE[31]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \Q[112]_i_1 
       (.I0(STALL_EN),
        .I1(\Q[112]_i_2_n_0 ),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[4]),
        .I5(EX_BR_TAKEN),
        .O(ID_EX_D[112]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'hFF02FFFF)) 
    \Q[112]_i_2 
       (.I0(I_MEM_DOUT_IBUF[13]),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[2]),
        .O(\Q[112]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFEFFFFF)) 
    \Q[113]_i_1 
       (.I0(I_MEM_DOUT_IBUF[3]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[5]),
        .I3(I_MEM_DOUT_IBUF[4]),
        .I4(\Q[125]_i_2_n_0 ),
        .I5(STALL_EN),
        .O(ID_WB_AFTER_LU));
  LUT6 #(
    .INIT(64'h8000800080808000)) 
    \Q[114]_i_1 
       (.I0(I_MEM_DOUT_IBUF[12]),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .I5(I_MEM_DOUT_IBUF[2]),
        .O(DECODED_INSTRUCTION[20]));
  LUT6 #(
    .INIT(64'h0000F40000000000)) 
    \Q[115]_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[4]),
        .I2(EX_BR_TAKEN),
        .I3(I_MEM_DOUT_IBUF[13]),
        .I4(I_MEM_DOUT_IBUF[12]),
        .I5(I_MEM_DOUT_IBUF[14]),
        .O(DECODED_INSTRUCTION[21]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT5 #(
    .INIT(32'h00004000)) 
    \Q[116]_i_1 
       (.I0(\Q[123]_i_3_n_0 ),
        .I1(I_MEM_DOUT_IBUF[14]),
        .I2(I_MEM_DOUT_IBUF[30]),
        .I3(I_MEM_DOUT_IBUF[12]),
        .I4(I_MEM_DOUT_IBUF[13]),
        .O(DECODED_INSTRUCTION[22]));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \Q[117]_i_1 
       (.I0(\Q[123]_i_3_n_0 ),
        .I1(I_MEM_DOUT_IBUF[14]),
        .I2(I_MEM_DOUT_IBUF[30]),
        .I3(I_MEM_DOUT_IBUF[12]),
        .I4(I_MEM_DOUT_IBUF[13]),
        .O(DECODED_INSTRUCTION[23]));
  LUT6 #(
    .INIT(64'h0000551000000000)) 
    \Q[118]_i_1 
       (.I0(I_MEM_DOUT_IBUF[13]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[4]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[12]),
        .I5(I_MEM_DOUT_IBUF[14]),
        .O(DECODED_INSTRUCTION[24]));
  LUT6 #(
    .INIT(64'h0800080008080800)) 
    \Q[119]_i_1 
       (.I0(I_MEM_DOUT_IBUF[12]),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .I5(I_MEM_DOUT_IBUF[2]),
        .O(DECODED_INSTRUCTION[25]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[11]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [11]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [10]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [11]));
  LUT6 #(
    .INIT(64'h000000008A888A8A)) 
    \Q[11]_i_10 
       (.I0(\Q[11]_i_16_n_0 ),
        .I1(\Q[67]_i_12_n_0 ),
        .I2(\Q[11]_i_17_n_0 ),
        .I3(\Q[21]_i_10__0_n_0 ),
        .I4(\Q[35]_i_32_n_0 ),
        .I5(\Q[29]_i_7_n_0 ),
        .O(\Q[11]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \Q[11]_i_11 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4447474774777777)) 
    \Q[11]_i_16 
       (.I0(\Q[35]_i_26_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[31]_i_13__0_n_0 ),
        .I4(\Q[35]_i_28_n_0 ),
        .I5(\Q[35]_i_29_n_0 ),
        .O(\Q[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB800B800B800)) 
    \Q[11]_i_17 
       (.I0(\custom_alu/int2fp/INT_VAL0 [4]),
        .I1(PSUM3__0_carry__0_i_10__2_n_0),
        .I2(ALU_DIN1[4]),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[31]_i_11__0_n_0 ),
        .O(\Q[11]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[11]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[12] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/data23 [11]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\Q[11]_i_2__0_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [11]));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \Q[11]_i_1__1 
       (.I0(\Q[11]_i_2_n_0 ),
        .I1(\Q[11]_i_3_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\Q[11]_i_4__0_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[6]),
        .O(data0[6]));
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \Q[11]_i_1__2 
       (.I0(\Q[11]_i_2__1_n_0 ),
        .I1(\Q[11]_i_3__0_n_0 ),
        .I2(\Q[11]_i_4__1_n_0 ),
        .I3(\Q[11]_i_5__1_n_0 ),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(EX_MEM_Q[11]),
        .O(data1[6]));
  LUT6 #(
    .INIT(64'h0D0D0D0D000D0D0D)) 
    \Q[11]_i_2 
       (.I0(\Q[14]_i_4__0_n_0 ),
        .I1(INT0_carry__0_i_8_n_0),
        .I2(\Q[11]_i_5__0_n_0 ),
        .I3(\Q[11]_i_6__0_n_0 ),
        .I4(\Q[27]_i_7_n_0 ),
        .I5(\Q[11]_i_7__0_n_0 ),
        .O(\Q[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBBB8B8B8)) 
    \Q[11]_i_2__0 
       (.I0(\custom_alu/fp32_add/sel0 [11]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\Q[11]_i_3__1_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [10]),
        .O(\Q[11]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[11]_i_2__1 
       (.I0(D_MEM_DOUT_IBUF[14]),
        .I1(D_MEM_DOUT_IBUF[6]),
        .I2(D_MEM_DOUT_IBUF[30]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[22]),
        .O(\Q[11]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[11]_i_3 
       (.I0(\custom_alu/fp32_mult/product_mantissa [6]),
        .I1(\Q[65]_i_5_n_0 ),
        .O(\Q[11]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'hDC)) 
    \Q[11]_i_3__0 
       (.I0(MEM_LOAD_SEL[5]),
        .I1(MEM_LOAD_SEL[6]),
        .I2(MEM_LOAD_SEL[2]),
        .O(\Q[11]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h5555510100005101)) 
    \Q[11]_i_3__1 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .I1(\Q[11]_i_4_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [8]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [9]),
        .O(\Q[11]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF7400000074)) 
    \Q[11]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\Q[11]_i_5_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [18]),
        .I4(\custom_alu/fp32_add/sel0 [19]),
        .I5(\Q[11]_i_6_n_0 ),
        .O(\Q[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB8B8888BB8B)) 
    \Q[11]_i_4__0 
       (.I0(\custom_alu/MULT [6]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(EX_CUSTOM_ALU_SEL[29]),
        .I3(\custom_alu/Q [6]),
        .I4(EX_CUSTOM_ALU_SEL[30]),
        .I5(\custom_alu/MULT [38]),
        .O(\Q[11]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[11]_i_4__1 
       (.I0(D_MEM_DOUT_IBUF[6]),
        .I1(D_MEM_DOUT_IBUF[22]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[30]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[14]),
        .O(\Q[11]_i_4__1_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[11]_i_5 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [16]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [15]),
        .I4(\Q[11]_i_7_n_0 ),
        .O(\Q[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[11]_i_5__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [6]),
        .O(\Q[11]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'h23)) 
    \Q[11]_i_5__1 
       (.I0(MEM_LOAD_SEL[5]),
        .I1(MEM_LOAD_SEL[6]),
        .I2(MEM_LOAD_SEL[2]),
        .O(\Q[11]_i_5__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \Q[11]_i_6 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [6]),
        .O(\Q[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h07070700FFFFFFFF)) 
    \Q[11]_i_6__0 
       (.I0(\Q[35]_i_21_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[11]_i_9_n_0 ),
        .I3(\Q[11]_i_10_n_0 ),
        .I4(\Q[11]_i_11_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[11]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h4444477777774777)) 
    \Q[11]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [14]),
        .I2(\custom_alu/fp32_add/sel0 [12]),
        .I3(\custom_alu/fp32_add/sel0 [0]),
        .I4(\custom_alu/fp32_add/sel0 [13]),
        .I5(\custom_alu/fp32_add/sel0 [1]),
        .O(\Q[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[11]_i_7__0 
       (.I0(\Q[28]_i_18_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_20_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[35]_i_19_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[11]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h0000CCA0)) 
    \Q[11]_i_9 
       (.I0(ALU_DIN1[0]),
        .I1(\Q[47]_i_9_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[27]_i_13_n_0 ),
        .O(\Q[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AE00)) 
    \Q[120]_i_1 
       (.I0(EX_BR_TAKEN),
        .I1(I_MEM_DOUT_IBUF[4]),
        .I2(I_MEM_DOUT_IBUF[2]),
        .I3(I_MEM_DOUT_IBUF[13]),
        .I4(I_MEM_DOUT_IBUF[12]),
        .I5(I_MEM_DOUT_IBUF[14]),
        .O(DECODED_INSTRUCTION[26]));
  LUT6 #(
    .INIT(64'h1000100010101000)) 
    \Q[121]_i_1 
       (.I0(I_MEM_DOUT_IBUF[14]),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[12]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .I5(I_MEM_DOUT_IBUF[2]),
        .O(DECODED_INSTRUCTION[27]));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \Q[122]_i_1 
       (.I0(\Q[123]_i_3_n_0 ),
        .I1(I_MEM_DOUT_FILTERED[5]),
        .I2(I_MEM_DOUT_IBUF[30]),
        .I3(I_MEM_DOUT_IBUF[13]),
        .I4(I_MEM_DOUT_IBUF[12]),
        .I5(I_MEM_DOUT_IBUF[14]),
        .O(DECODED_INSTRUCTION[28]));
  LUT6 #(
    .INIT(64'hAFBFAFAFABBBAAAA)) 
    \Q[123]_i_1 
       (.I0(ID_MEM),
        .I1(\Q[123]_i_3_n_0 ),
        .I2(I_MEM_DOUT_FILTERED[5]),
        .I3(I_MEM_DOUT_IBUF[30]),
        .I4(\Q[123]_i_5_n_0 ),
        .I5(\Q[123]_i_6_n_0 ),
        .O(DECODED_INSTRUCTION[29]));
  LUT6 #(
    .INIT(64'h0000000100000101)) 
    \Q[123]_i_2 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[3]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[2]),
        .I4(EX_BR_TAKEN),
        .I5(\Q[160]_i_2_n_0 ),
        .O(ID_MEM));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'h0B)) 
    \Q[123]_i_3 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[4]),
        .I2(EX_BR_TAKEN),
        .O(\Q[123]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \Q[123]_i_4 
       (.I0(EX_BR_TAKEN),
        .I1(I_MEM_DOUT_IBUF[5]),
        .O(I_MEM_DOUT_FILTERED[5]));
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \Q[123]_i_5 
       (.I0(I_MEM_DOUT_IBUF[14]),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[13]),
        .O(\Q[123]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \Q[123]_i_6 
       (.I0(I_MEM_DOUT_IBUF[3]),
        .I1(I_MEM_DOUT_IBUF[6]),
        .I2(I_MEM_DOUT_IBUF[2]),
        .I3(I_MEM_DOUT_IBUF[4]),
        .I4(EX_BR_TAKEN),
        .O(\Q[123]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hF6)) 
    \Q[124]_i_1 
       (.I0(ID_WE_AFTER_LU3),
        .I1(STALL_EN),
        .I2(\Q[124]_i_3_n_0 ),
        .O(ID_EX_D[124]));
  LUT6 #(
    .INIT(64'h0000000000010501)) 
    \Q[124]_i_2 
       (.I0(\Q[161]_i_4_n_0 ),
        .I1(I_MEM_DOUT_FILTERED[2]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .I3(I_MEM_DOUT_IBUF[13]),
        .I4(I_MEM_DOUT_IBUF[12]),
        .I5(\Q[161]_i_2_n_0 ),
        .O(ID_WE_AFTER_LU3));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    \Q[124]_i_3 
       (.I0(LU_HAZARD),
        .I1(\Q[112]_i_2_n_0 ),
        .I2(EX_BR_TAKEN),
        .I3(I_MEM_DOUT_IBUF[5]),
        .I4(I_MEM_DOUT_IBUF[4]),
        .I5(\Q[161]_i_2_n_0 ),
        .O(\Q[124]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5155515100000000)) 
    \Q[125]_i_1 
       (.I0(STALL_EN),
        .I1(\Q[125]_i_2_n_0 ),
        .I2(\Q[161]_i_4_n_0 ),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[3]),
        .I5(ID_BR),
        .O(ID_JAL_AFTER_LU));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \Q[125]_i_2 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[6]),
        .O(\Q[125]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT5 #(
    .INIT(32'hFFFFFFA2)) 
    \Q[125]_i_3 
       (.I0(\Q[90]_i_4_n_0 ),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .I3(DECODED_INSTRUCTION[13]),
        .I4(DECODED_INSTRUCTION[12]),
        .O(ID_BR));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \Q[125]_i_4 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[3]),
        .I3(I_MEM_DOUT_IBUF[6]),
        .I4(EX_BR_TAKEN),
        .I5(I_MEM_DOUT_IBUF[2]),
        .O(DECODED_INSTRUCTION[13]));
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[12]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [12]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [11]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [12]));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000008B)) 
    \Q[12]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [3]),
        .I1(\custom_alu/fp32_add/sel0 [14]),
        .I2(\Q[12]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [15]),
        .I4(\custom_alu/fp32_add/sel0 [16]),
        .I5(\Q[12]_i_13__0_n_0 ),
        .O(\Q[12]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[12]_i_11 
       (.I0(\Q[16]_i_16_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[12]_i_15_n_0 ),
        .O(\Q[12]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \Q[12]_i_11__0 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [7]),
        .O(\Q[12]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h0101000155555555)) 
    \Q[12]_i_11__1 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[67]_i_12_n_0 ),
        .I2(\Q[12]_i_18__0_n_0 ),
        .I3(\Q[29]_i_18__0_n_0 ),
        .I4(\Q[21]_i_10__0_n_0 ),
        .I5(\Q[12]_i_19__0_n_0 ),
        .O(\Q[12]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'h4744477747774777)) 
    \Q[12]_i_12 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [13]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [12]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .I5(\custom_alu/fp32_add/sel0 [0]),
        .O(\Q[12]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFB8880000B888)) 
    \Q[12]_i_12__0 
       (.I0(\Q[47]_i_9_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[17]_i_10__0_n_0 ),
        .I3(ALU_DIN1[0]),
        .I4(\Q[28]_i_11_n_0 ),
        .I5(\Q[35]_i_32_n_0 ),
        .O(\Q[12]_i_12__0_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \Q[12]_i_12__1 
       (.I0(\Q[16]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[12]_i_16_n_0 ),
        .I3(\Q[16]_i_20_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[12]_i_12__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[12]_i_13 
       (.I0(\Q[16]_i_19_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[12]_i_17_n_0 ),
        .O(\Q[12]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF088)) 
    \Q[12]_i_13__0 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [5]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[12]_i_13__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000777)) 
    \Q[12]_i_13__1 
       (.I0(\Q[28]_i_7_n_0 ),
        .I1(\Q[35]_i_20_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[28]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .O(\Q[12]_i_13__1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[12]_i_14 
       (.I0(\Q_reg[16]_i_13_n_7 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_18_n_4 ),
        .O(\Q[12]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \Q[12]_i_14__0 
       (.I0(\Q[12]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[12]_i_19_n_0 ),
        .I3(\Q[16]_i_18_n_0 ),
        .I4(\Q[12]_i_16_n_0 ),
        .I5(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[12]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[12]_i_15 
       (.I0(ALU_DIN2[19]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[19]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[12]_i_20_n_0 ),
        .O(\Q[12]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[12]_i_15__0 
       (.I0(\Q_reg[49]_i_18_n_4 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_18_n_5 ),
        .O(\Q[12]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[12]_i_16 
       (.I0(ALU_DIN2[18]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[18]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[4]_i_24_n_0 ),
        .O(\Q[12]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[12]_i_16__0 
       (.I0(\Q_reg[49]_i_18_n_5 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_18_n_6 ),
        .O(\Q[12]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[12]_i_17 
       (.I0(ALU_DIN2[17]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[17]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[12]_i_21_n_0 ),
        .O(\Q[12]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[12]_i_17__0 
       (.I0(\Q_reg[49]_i_18_n_6 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_18_n_7 ),
        .O(\Q[12]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[12]_i_18 
       (.I0(ALU_DIN2[20]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[20]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[12]_i_22_n_0 ),
        .O(\Q[12]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \Q[12]_i_18__0 
       (.I0(\Q[35]_i_28_n_0 ),
        .I1(\Q[31]_i_14__0_n_0 ),
        .I2(ALU_DIN1[4]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [4]),
        .I5(\Q[31]_i_11__0_n_0 ),
        .O(\Q[12]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[12]_i_19 
       (.I0(ALU_DIN2[16]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[16]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[4]_i_22_n_0 ),
        .O(\Q[12]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFD0D0000FD0D)) 
    \Q[12]_i_19__0 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[35]_i_27_n_0 ),
        .O(\Q[12]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[12]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[13] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/data23 [12]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\Q[12]_i_3__0_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [12]));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \Q[12]_i_1__1 
       (.I0(\Q[12]_i_2_n_0 ),
        .I1(\Q[12]_i_3__1_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\Q[12]_i_4__1_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[7]),
        .O(data0[7]));
  LUT4 #(
    .INIT(16'hFB08)) 
    \Q[12]_i_1__2 
       (.I0(\Q[12]_i_2__0_n_0 ),
        .I1(EX_MEM_Q[39]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[12]),
        .O(data1[7]));
  LUT6 #(
    .INIT(64'h2222222220200020)) 
    \Q[12]_i_2 
       (.I0(\Q[12]_i_5__2_n_0 ),
        .I1(\Q[12]_i_6__1_n_0 ),
        .I2(\Q[26]_i_7_n_0 ),
        .I3(\Q[12]_i_7__0_n_0 ),
        .I4(\Q[12]_i_8_n_0 ),
        .I5(\Q[12]_i_9__0_n_0 ),
        .O(\Q[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[12]_i_20 
       (.I0(EX_RF_RD2[11]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[90]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[11]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[12]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[12]_i_21 
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[88]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[9]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[12]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[12]_i_22 
       (.I0(EX_RF_RD2[12]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[91]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[12]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[12]_i_22_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT5 #(
    .INIT(32'hCCAACCCA)) 
    \Q[12]_i_2__0 
       (.I0(\Q[12]_i_3__2_n_0 ),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(MEM_LOAD_SEL[2]),
        .I3(MEM_LOAD_SEL[6]),
        .I4(MEM_LOAD_SEL[5]),
        .O(\Q[12]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[12]_i_2__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[12]),
        .I2(STALL_EN),
        .I3(IF_PC2[12]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[12] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[12]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[12]_i_3 
       (.I0(\Q[12]_i_11_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\Q[16]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[16]_i_15__0_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [11]));
  LUT5 #(
    .INIT(32'hBBB8B8B8)) 
    \Q[12]_i_3__0 
       (.I0(\custom_alu/fp32_add/sel0 [12]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\Q[12]_i_8__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[12]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[12]_i_3__1 
       (.I0(\custom_alu/fp32_mult/product_mantissa [7]),
        .I1(\Q[65]_i_5_n_0 ),
        .O(\Q[12]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[12]_i_3__2 
       (.I0(D_MEM_DOUT_IBUF[7]),
        .I1(D_MEM_DOUT_IBUF[23]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[31]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[15]),
        .O(\Q[12]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[12]_i_3__3 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[11]),
        .I2(STALL_EN),
        .I3(IF_PC2[11]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[11] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[12]_i_3__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[12]_i_4 
       (.I0(\Q[12]_i_12__1_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[12]_i_11_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[16]_i_14_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [10]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[12]_i_4__0 
       (.I0(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[12]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB8B8888BB8B)) 
    \Q[12]_i_4__1 
       (.I0(\custom_alu/MULT [7]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(EX_CUSTOM_ALU_SEL[29]),
        .I3(\custom_alu/Q [7]),
        .I4(EX_CUSTOM_ALU_SEL[30]),
        .I5(\custom_alu/MULT [39]),
        .O(\Q[12]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[12]_i_4__2 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[10]),
        .I2(STALL_EN),
        .I3(IF_PC2[10]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[10] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[12]_i_4__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[12]_i_5 
       (.I0(\Q[12]_i_13_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\Q[12]_i_11_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[12]_i_12__1_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [9]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[12]_i_5__0 
       (.I0(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[12]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[12]_i_5__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[9]),
        .I2(STALL_EN),
        .I3(IF_PC2[9]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[9] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[12]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0047FFFFFFFF)) 
    \Q[12]_i_5__2 
       (.I0(INT0_carry__0_i_5_n_0),
        .I1(ALU_DIN1[23]),
        .I2(INT0_carry__0_i_7_n_0),
        .I3(INT0_carry_i_6_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[12]_i_5__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[12]_i_6 
       (.I0(\Q[12]_i_14__0_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[12]_i_13_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[12]_i_11_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [8]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[12]_i_6__0 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .O(\Q[12]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[12]_i_6__1 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [7]),
        .O(\Q[12]_i_6__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[12]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [9]),
        .O(\Q[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEEFFFFEFEE)) 
    \Q[12]_i_7__0 
       (.I0(\Q[12]_i_11__1_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[35]_i_21_n_0 ),
        .I3(\Q[28]_i_12_n_0 ),
        .I4(\Q[28]_i_21_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[12]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h888F8888)) 
    \Q[12]_i_8 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[27]_i_13_n_0 ),
        .I3(\Q[22]_i_7__0_n_0 ),
        .I4(\Q[12]_i_12__0_n_0 ),
        .O(\Q[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5555510100005101)) 
    \Q[12]_i_8__0 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .I1(\Q[12]_i_9_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [9]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [10]),
        .O(\Q[12]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF4F0000004F)) 
    \Q[12]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\Q[12]_i_10_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [18]),
        .I4(\custom_alu/fp32_add/sel0 [19]),
        .I5(\Q[12]_i_11__0_n_0 ),
        .O(\Q[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF4540FFFFFFFF)) 
    \Q[12]_i_9__0 
       (.I0(\Q[12]_i_13__1_n_0 ),
        .I1(\Q[17]_i_11__0_n_0 ),
        .I2(\Q[28]_i_6_n_0 ),
        .I3(\Q[26]_i_15__0_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[12]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[13]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [13]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [12]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [13]));
  LUT6 #(
    .INIT(64'h000000008A888A8A)) 
    \Q[13]_i_10 
       (.I0(\Q[13]_i_15_n_0 ),
        .I1(\Q[67]_i_12_n_0 ),
        .I2(\Q[13]_i_16_n_0 ),
        .I3(\Q[21]_i_10__0_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .I5(\Q[29]_i_7_n_0 ),
        .O(\Q[13]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \Q[13]_i_11 
       (.I0(\Q[27]_i_13_n_0 ),
        .I1(\Q[69]_i_20_n_0 ),
        .O(\Q[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \Q[13]_i_12 
       (.I0(ALU_DIN1[0]),
        .I1(EX_RF_RD1[15]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[141]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\custom_alu/int2fp/INT_VAL0 [15]),
        .O(\Q[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFB00FBFF0B000B)) 
    \Q[13]_i_13 
       (.I0(\Q[47]_i_9_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[35]_i_32_n_0 ),
        .O(\Q[13]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00000777)) 
    \Q[13]_i_14 
       (.I0(\Q[28]_i_7_n_0 ),
        .I1(\Q[28]_i_18_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[17]_i_11__0_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .O(\Q[13]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4447474774777777)) 
    \Q[13]_i_15 
       (.I0(\Q[35]_i_22_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[31]_i_13__0_n_0 ),
        .I4(\Q[35]_i_26_n_0 ),
        .I5(\Q[35]_i_27_n_0 ),
        .O(\Q[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \Q[13]_i_16 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[31]_i_14__0_n_0 ),
        .I2(ALU_DIN1[5]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [5]),
        .I5(\Q[31]_i_11__0_n_0 ),
        .O(\Q[13]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000EEF0)) 
    \Q[13]_i_1__0 
       (.I0(\Q[13]_i_2_n_0 ),
        .I1(\Q[13]_i_3__0_n_0 ),
        .I2(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[14] ),
        .I3(\Q[30]_i_2__1_n_0 ),
        .I4(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [13]));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \Q[13]_i_1__1 
       (.I0(\Q[13]_i_2__0_n_0 ),
        .I1(\Q[13]_i_3_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\Q[13]_i_4_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[8]),
        .O(data0[8]));
  LUT6 #(
    .INIT(64'hFFFFF8FF0000F800)) 
    \Q[13]_i_1__2 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(\Q[13]_i_2__1_n_0 ),
        .I3(EX_MEM_Q[39]),
        .I4(EX_MEM_Q[37]),
        .I5(EX_MEM_Q[13]),
        .O(data1[8]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[13]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [13]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [13]),
        .O(\Q[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h2222222220200020)) 
    \Q[13]_i_2__0 
       (.I0(\Q[13]_i_5__0_n_0 ),
        .I1(\Q[13]_i_6__0_n_0 ),
        .I2(\Q[26]_i_7_n_0 ),
        .I3(\Q[13]_i_7__0_n_0 ),
        .I4(\Q[13]_i_8__0_n_0 ),
        .I5(\Q[13]_i_9__0_n_0 ),
        .O(\Q[13]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AA8080000A808)) 
    \Q[13]_i_2__1 
       (.I0(\Q[11]_i_5__1_n_0 ),
        .I1(D_MEM_DOUT_IBUF[8]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I3(D_MEM_DOUT_IBUF[24]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[16]),
        .O(\Q[13]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[13]_i_3 
       (.I0(\custom_alu/fp32_mult/product_mantissa [8]),
        .I1(\Q[65]_i_5_n_0 ),
        .O(\Q[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00F80000)) 
    \Q[13]_i_3__0 
       (.I0(\custom_alu/fp32_add/sel0 [12]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\Q[13]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [23]),
        .I4(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[13]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB8B8888BB8B)) 
    \Q[13]_i_4 
       (.I0(\custom_alu/MULT [8]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(EX_CUSTOM_ALU_SEL[29]),
        .I3(\custom_alu/Q [8]),
        .I4(EX_CUSTOM_ALU_SEL[30]),
        .I5(\custom_alu/MULT [40]),
        .O(\Q[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5555510100005101)) 
    \Q[13]_i_4__0 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .I1(\Q[13]_i_5_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [10]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[13]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'h02F20EFE)) 
    \Q[13]_i_5 
       (.I0(\Q[13]_i_6_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [19]),
        .I3(\custom_alu/fp32_add/sel0 [9]),
        .I4(\custom_alu/fp32_add/sel0 [8]),
        .O(\Q[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0047FFFFFFFF)) 
    \Q[13]_i_5__0 
       (.I0(INT0_carry__0_i_6_n_0),
        .I1(ALU_DIN1[23]),
        .I2(INT0_carry__0_i_5_n_0),
        .I3(INT0_carry_i_6_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[13]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4F4F4F4F44)) 
    \Q[13]_i_6 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\Q[13]_i_7_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\Q[13]_i_8_n_0 ),
        .O(\Q[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[13]_i_6__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [8]),
        .O(\Q[13]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF088)) 
    \Q[13]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [6]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEEFFFFEFEE)) 
    \Q[13]_i_7__0 
       (.I0(\Q[13]_i_10_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[35]_i_19_n_0 ),
        .I3(\Q[28]_i_12_n_0 ),
        .I4(\Q[28]_i_21_n_0 ),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[13]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[13]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [14]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [13]),
        .I4(\Q[13]_i_9_n_0 ),
        .O(\Q[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h888F8F8F88888888)) 
    \Q[13]_i_8__0 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[13]_i_11_n_0 ),
        .I3(\Q[13]_i_12_n_0 ),
        .I4(\Q[22]_i_7__0_n_0 ),
        .I5(\Q[13]_i_13_n_0 ),
        .O(\Q[13]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h4744477747774777)) 
    \Q[13]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [11]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [10]),
        .O(\Q[13]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF4540FFFFFFFF)) 
    \Q[13]_i_9__0 
       (.I0(\Q[13]_i_14_n_0 ),
        .I1(\Q[17]_i_14_n_0 ),
        .I2(\Q[28]_i_6_n_0 ),
        .I3(\Q[26]_i_15__0_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[13]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[14]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [14]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [13]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [14]));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[14]_i_1__0 
       (.I0(\Q[14]_i_2_n_0 ),
        .I1(\Q[14]_i_3_n_0 ),
        .I2(\Q[14]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[15] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [14]));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[14]_i_1__1 
       (.I0(\Q[14]_i_2__0_n_0 ),
        .I1(\Q[14]_i_3__0_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[9]),
        .O(data0[9]));
  LUT6 #(
    .INIT(64'hFFFFF8FF0000F800)) 
    \Q[14]_i_1__2 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(\Q[14]_i_2__1_n_0 ),
        .I3(EX_MEM_Q[39]),
        .I4(EX_MEM_Q[37]),
        .I5(EX_MEM_Q[14]),
        .O(data1[9]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[14]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [14]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [14]),
        .O(\Q[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[14]_i_2__0 
       (.I0(\custom_alu/MULT [9]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [41]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [9]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[14]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AA8080000A808)) 
    \Q[14]_i_2__1 
       (.I0(\Q[11]_i_5__1_n_0 ),
        .I1(D_MEM_DOUT_IBUF[9]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I3(D_MEM_DOUT_IBUF[25]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[17]),
        .O(\Q[14]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFFCDDFCCCFCDD)) 
    \Q[14]_i_3 
       (.I0(\Q[14]_i_5_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [12]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hDDD0DDDDDDD0DDD0)) 
    \Q[14]_i_3__0 
       (.I0(\custom_alu/fp32_mult/product_mantissa [9]),
        .I1(\Q[65]_i_5_n_0 ),
        .I2(\Q[24]_i_6__0_n_0 ),
        .I3(\Q[24]_i_7__0_n_0 ),
        .I4(INT0_carry__1_i_9_n_0),
        .I5(\Q[14]_i_4__0_n_0 ),
        .O(\Q[14]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT4 #(
    .INIT(16'hF4FF)) 
    \Q[14]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [13]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [23]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[14]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT4 #(
    .INIT(16'h02A2)) 
    \Q[14]_i_4__0 
       (.I0(EX_CUSTOM_ALU_SEL[27]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .O(\Q[14]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'h02F20EFE)) 
    \Q[14]_i_5 
       (.I0(\Q[14]_i_6_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [19]),
        .I3(\custom_alu/fp32_add/sel0 [10]),
        .I4(\custom_alu/fp32_add/sel0 [9]),
        .O(\Q[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[14]_i_6 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [7]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\Q[14]_i_7_n_0 ),
        .O(\Q[14]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[14]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [5]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\Q[14]_i_8_n_0 ),
        .O(\Q[14]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[14]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [13]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [12]),
        .I4(\Q[14]_i_9_n_0 ),
        .O(\Q[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4744477747774777)) 
    \Q[14]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [11]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [10]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [9]),
        .O(\Q[14]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT5 #(
    .INIT(32'h00AB00AF)) 
    \Q[158]_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .O(ID_IMMEDIATE_EN));
  LUT5 #(
    .INIT(32'h00AB00AF)) 
    \Q[158]_rep__0_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .O(\Q[158]_rep__0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00AB00AF)) 
    \Q[158]_rep__1_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .O(\Q[158]_rep__1_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00AB00AF)) 
    \Q[158]_rep__2_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .O(\Q[158]_rep__2_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00AB00AF)) 
    \Q[158]_rep__3_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .O(\Q[158]_rep__3_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00AB00AF)) 
    \Q[158]_rep__4_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .O(\Q[158]_rep__4_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00AB00AF)) 
    \Q[158]_rep_i_1 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[4]),
        .O(\Q[158]_rep_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[15]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [15]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [14]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [15]));
  LUT6 #(
    .INIT(64'h4744477747774777)) 
    \Q[15]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [10]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [9]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [8]),
        .O(\Q[15]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5400)) 
    \Q[15]_i_12 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[15]_i_17_n_0 ),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[15]_i_18_n_0 ),
        .I4(\Q[15]_i_19_n_0 ),
        .O(\Q[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B0B0)) 
    \Q[15]_i_13 
       (.I0(\Q[29]_i_18__0_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[15]_i_20_n_0 ),
        .I3(\Q[17]_i_15_n_0 ),
        .I4(\Q[69]_i_16_n_0 ),
        .I5(\Q[28]_i_11_n_0 ),
        .O(\Q[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFFFEEEEEEEE)) 
    \Q[15]_i_14 
       (.I0(\Q[69]_i_20_n_0 ),
        .I1(\Q[27]_i_13_n_0 ),
        .I2(\custom_alu/int2fp/INT_VAL0 [5]),
        .I3(ALU_DIN1[31]),
        .I4(ALU_DIN1[5]),
        .I5(\Q[28]_i_11_n_0 ),
        .O(\Q[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \Q[15]_i_15 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(EX_RF_RD1[14]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[140]),
        .I4(ALU_DIN1[31]),
        .I5(\custom_alu/int2fp/INT_VAL0 [14]),
        .O(\Q[15]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[15]_i_16 
       (.I0(\Q[69]_i_16_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[17]_i_10__0_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[15]_i_17 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[35]_i_27_n_0 ),
        .O(\Q[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h4447474774777777)) 
    \Q[15]_i_18 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[31]_i_13__0_n_0 ),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[15]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \Q[15]_i_19 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[28]_i_18_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[15]_i_1__0 
       (.I0(\Q[15]_i_2_n_0 ),
        .I1(\Q[15]_i_3_n_0 ),
        .I2(\Q[15]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[16] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[15]_i_1__1 
       (.I0(\Q[15]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[0]),
        .I5(\Q[15]_i_3__1_n_0 ),
        .O(ID_RD2_FORWARDED[0]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[15]_i_1__2 
       (.I0(\Q[15]_i_2__0_n_0 ),
        .I1(\Q[15]_i_3__0_n_0 ),
        .I2(\Q[15]_i_4__0_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[10]),
        .O(data0[10]));
  LUT6 #(
    .INIT(64'hFFFFF8FF0000F800)) 
    \Q[15]_i_1__3 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(\Q[15]_i_2__2_n_0 ),
        .I3(EX_MEM_Q[39]),
        .I4(EX_MEM_Q[37]),
        .I5(EX_MEM_Q[15]),
        .O(data1[10]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[15]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [15]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [15]),
        .O(\Q[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00E0E0)) 
    \Q[15]_i_20 
       (.I0(\Q[28]_i_18_n_0 ),
        .I1(\Q[17]_i_11__0_n_0 ),
        .I2(\Q[15]_i_21_n_0 ),
        .I3(\Q[35]_i_32_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[17]_i_10__0_n_0 ),
        .O(\Q[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAFCCAFFFA0CCA000)) 
    \Q[15]_i_21 
       (.I0(\custom_alu/int2fp/INT_VAL0 [1]),
        .I1(ALU_DIN1[1]),
        .I2(\custom_alu/int2fp/INT_VAL0 [14]),
        .I3(ALU_DIN1[31]),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN1[0]),
        .O(\Q[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[15]_i_2__0 
       (.I0(\custom_alu/MULT [10]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [42]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [10]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[15]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[15]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[0]),
        .I2(CRF_RD2_IBUF[0]),
        .I3(RF_RD2_IBUF[0]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[15]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AA8080000A808)) 
    \Q[15]_i_2__2 
       (.I0(\Q[11]_i_5__1_n_0 ),
        .I1(D_MEM_DOUT_IBUF[10]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I3(D_MEM_DOUT_IBUF[26]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[18]),
        .O(\Q[15]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFFCDDFCCCFCDD)) 
    \Q[15]_i_3 
       (.I0(\Q[15]_i_5_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [13]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[15]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \Q[15]_i_3__0 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [10]),
        .O(\Q[15]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[15]_i_3__1 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(data1[0]),
        .O(\Q[15]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT4 #(
    .INIT(16'hF4FF)) 
    \Q[15]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [14]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [23]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0E000E0F0E000E00)) 
    \Q[15]_i_4__0 
       (.I0(ALU_DIN1[31]),
        .I1(INT0_carry__1_i_8_n_0),
        .I2(\Q[15]_i_6__0_n_0 ),
        .I3(EX_CUSTOM_ALU_SEL[27]),
        .I4(\Q[15]_i_7__0_n_0 ),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[15]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'h02F20EFE)) 
    \Q[15]_i_5 
       (.I0(\Q[15]_i_6_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [19]),
        .I3(\custom_alu/fp32_add/sel0 [11]),
        .I4(\custom_alu/fp32_add/sel0 [10]),
        .O(\Q[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h5554FFFF55545554)) 
    \Q[15]_i_6 
       (.I0(\Q[15]_i_7_n_0 ),
        .I1(\Q[15]_i_8_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [16]),
        .I3(\custom_alu/fp32_add/sel0 [15]),
        .I4(\custom_alu/fp32_add/sel0 [9]),
        .I5(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[15]_i_6__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [10]),
        .O(\Q[15]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF088)) 
    \Q[15]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [8]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555DD5D)) 
    \Q[15]_i_7__0 
       (.I0(\Q[26]_i_7_n_0 ),
        .I1(\Q[15]_i_12_n_0 ),
        .I2(\Q[15]_i_13_n_0 ),
        .I3(\Q[15]_i_14_n_0 ),
        .I4(\Q[15]_i_15_n_0 ),
        .I5(\Q[15]_i_16_n_0 ),
        .O(\Q[15]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[15]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [14]),
        .I2(\custom_alu/fp32_add/sel0 [5]),
        .I3(\custom_alu/fp32_add/sel0 [13]),
        .I4(\Q[15]_i_9_n_0 ),
        .O(\Q[15]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[15]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [11]),
        .I4(\Q[15]_i_10_n_0 ),
        .O(\Q[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \Q[160]_i_1 
       (.I0(I_MEM_DOUT_IBUF[3]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[4]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(\Q[160]_i_2_n_0 ),
        .O(DECODED_INSTRUCTION[2]));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \Q[160]_i_2 
       (.I0(I_MEM_DOUT_IBUF[14]),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[13]),
        .O(\Q[160]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \Q[161]_i_1 
       (.I0(\Q[161]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[13]),
        .I3(I_MEM_DOUT_IBUF[14]),
        .I4(I_MEM_DOUT_FILTERED[2]),
        .I5(\Q[161]_i_4_n_0 ),
        .O(DECODED_INSTRUCTION[3]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \Q[161]_i_2 
       (.I0(I_MEM_DOUT_IBUF[3]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[6]),
        .O(\Q[161]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[161]_i_3 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[2]));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \Q[161]_i_4 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(EX_BR_TAKEN),
        .O(\Q[161]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \Q[164]_i_1 
       (.I0(I_MEM_DOUT_IBUF[12]),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[5]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[14]),
        .I5(\Q[169]_i_2_n_0 ),
        .O(DECODED_INSTRUCTION[6]));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \Q[165]_i_1 
       (.I0(I_MEM_DOUT_IBUF[14]),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[5]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[13]),
        .I5(\Q[169]_i_2_n_0 ),
        .O(DECODED_INSTRUCTION[7]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \Q[168]_i_1 
       (.I0(I_MEM_DOUT_IBUF[14]),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[13]),
        .I3(I_MEM_DOUT_IBUF[5]),
        .I4(EX_BR_TAKEN),
        .I5(\Q[169]_i_2_n_0 ),
        .O(DECODED_INSTRUCTION[10]));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \Q[169]_i_1 
       (.I0(EX_BR_TAKEN),
        .I1(I_MEM_DOUT_IBUF[5]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .I3(I_MEM_DOUT_IBUF[12]),
        .I4(I_MEM_DOUT_IBUF[13]),
        .I5(\Q[169]_i_2_n_0 ),
        .O(DECODED_INSTRUCTION[11]));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \Q[169]_i_2 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[3]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[2]),
        .O(\Q[169]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[16]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [16]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [15]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [16]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[16]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [13]),
        .O(\Q[16]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[16]_i_10__0 
       (.I0(\Q_reg[16]_i_13_n_4 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[16]_i_13_n_5 ),
        .O(\Q[16]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \Q[16]_i_11 
       (.I0(\Q[20]_i_19_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[16]_i_16_n_0 ),
        .O(\Q[16]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4F4F4F4F44)) 
    \Q[16]_i_11__0 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\Q[16]_i_12__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\Q[16]_i_13_n_0 ),
        .O(\Q[16]_i_11__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[16]_i_11__1 
       (.I0(\Q_reg[16]_i_13_n_5 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[16]_i_13_n_6 ),
        .O(\Q[16]_i_11__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[16]_i_12 
       (.I0(\Q[23]_i_19_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[16]_i_17_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [3]),
        .O(\Q[16]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF088)) 
    \Q[16]_i_12__0 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [9]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[16]_i_12__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[16]_i_12__1 
       (.I0(\Q_reg[16]_i_13_n_6 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[16]_i_13_n_7 ),
        .O(\Q[16]_i_12__1_n_0 ));
  LUT6 #(
    .INIT(64'h55305530553F5530)) 
    \Q[16]_i_13 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [6]),
        .I2(\custom_alu/fp32_add/sel0 [13]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\Q[16]_i_14__0_n_0 ),
        .I5(\Q[16]_i_15_n_0 ),
        .O(\Q[16]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00002F202F20)) 
    \Q[16]_i_13__0 
       (.I0(\Q[20]_i_20_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[16]_i_18_n_0 ),
        .I4(\Q[20]_i_21_n_0 ),
        .I5(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[16]_i_13__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \Q[16]_i_14 
       (.I0(\Q[16]_i_17_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[16]_i_19_n_0 ),
        .O(\Q[16]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \Q[16]_i_14__0 
       (.I0(\custom_alu/fp32_add/sel0 [12]),
        .I1(\Q[16]_i_16__0_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [10]),
        .I3(\custom_alu/fp32_add/sel0 [3]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .I5(\custom_alu/fp32_add/sel0 [4]),
        .O(\Q[16]_i_14__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[16]_i_15 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[16]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \Q[16]_i_15__0 
       (.I0(\Q[20]_i_20_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[16]_i_18_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I5(\Q[16]_i_20_n_0 ),
        .O(\Q[16]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h88888888BBB888B8)) 
    \Q[16]_i_16 
       (.I0(\Q[23]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(ALU_DIN2[15]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[15]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[16]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[16]_i_16__0 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [9]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [8]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [7]),
        .O(\Q[16]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[16]_i_17 
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[96]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[17]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[16]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[16]_i_18 
       (.I0(ALU_DIN2[22]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[22]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[16]_i_21_n_0 ),
        .O(\Q[16]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[16]_i_19 
       (.I0(ALU_DIN2[21]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[21]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[16]_i_22_n_0 ),
        .O(\Q[16]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[16]_i_1__0 
       (.I0(\Q[16]_i_2_n_0 ),
        .I1(\Q[16]_i_3__0_n_0 ),
        .I2(\Q[16]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[17] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [16]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[16]_i_1__1 
       (.I0(\Q[16]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[1]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[1]),
        .I5(\Q[16]_i_3__2_n_0 ),
        .O(ID_RD2_FORWARDED[1]));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[16]_i_1__2 
       (.I0(\Q[16]_i_2__0_n_0 ),
        .I1(\Q[16]_i_3__1_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[11]),
        .O(data0[11]));
  LUT6 #(
    .INIT(64'hFFFFF8FF0000F800)) 
    \Q[16]_i_1__3 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(\Q[16]_i_2__2_n_0 ),
        .I3(EX_MEM_Q[39]),
        .I4(EX_MEM_Q[37]),
        .I5(EX_MEM_Q[16]),
        .O(data1[11]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[16]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [16]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [16]),
        .O(\Q[16]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \Q[16]_i_20 
       (.I0(\Q[20]_i_22_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[12]_i_18_n_0 ),
        .O(\Q[16]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[16]_i_21 
       (.I0(EX_RF_RD2[14]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[93]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[14]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[16]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[16]_i_22 
       (.I0(EX_RF_RD2[13]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[92]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[13]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[16]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[16]_i_2__0 
       (.I0(\custom_alu/MULT [11]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [43]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(\custom_alu/Q [11]),
        .O(\Q[16]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[16]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[1]),
        .I2(CRF_RD2_IBUF[1]),
        .I3(RF_RD2_IBUF[1]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[16]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AA8080000A808)) 
    \Q[16]_i_2__2 
       (.I0(\Q[11]_i_5__1_n_0 ),
        .I1(D_MEM_DOUT_IBUF[11]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I3(D_MEM_DOUT_IBUF[27]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[19]),
        .O(\Q[16]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[16]_i_2__3 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[16]),
        .I2(STALL_EN),
        .I3(IF_PC2[16]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[16] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[16]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[16]_i_3 
       (.I0(\Q[16]_i_11_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\Q[16]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_14__1_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [15]));
  LUT6 #(
    .INIT(64'hFCFFFCDDFCCCFCDD)) 
    \Q[16]_i_3__0 
       (.I0(\Q[16]_i_6__0_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [14]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [13]),
        .O(\Q[16]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFF020000FF02FF02)) 
    \Q[16]_i_3__1 
       (.I0(\Q[26]_i_5__0_n_0 ),
        .I1(\Q[16]_i_4__1_n_0 ),
        .I2(\Q[16]_i_5__0_n_0 ),
        .I3(EX_CUSTOM_ALU_SEL[28]),
        .I4(\Q[65]_i_5_n_0 ),
        .I5(\custom_alu/fp32_mult/product_mantissa [11]),
        .O(\Q[16]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[16]_i_3__2 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(data1[1]),
        .O(\Q[16]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[16]_i_3__3 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[15]),
        .I2(STALL_EN),
        .I3(IF_PC2[15]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[15] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[16]_i_3__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[16]_i_4 
       (.I0(\Q[16]_i_13__0_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[16]_i_11_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[16]_i_12_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [14]));
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT4 #(
    .INIT(16'hF4FF)) 
    \Q[16]_i_4__0 
       (.I0(\custom_alu/fp32_add/sel0 [15]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [23]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[16]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'h80888000)) 
    \Q[16]_i_4__1 
       (.I0(\custom_alu/fp2int/INT0 [11]),
        .I1(EX_CUSTOM_ALU_SEL[27]),
        .I2(ID_EX_Q[157]),
        .I3(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I4(EX_RF_RD1[31]),
        .O(\Q[16]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[16]_i_4__2 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[14]),
        .I2(STALL_EN),
        .I3(IF_PC2[14]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[14] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[16]_i_4__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[16]_i_5 
       (.I0(\Q[16]_i_14_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\Q[16]_i_11_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[16]_i_13__0_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [13]));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \Q[16]_i_5__0 
       (.I0(\Q[27]_i_7_n_0 ),
        .I1(\Q[26]_i_11__0_n_0 ),
        .I2(\Q[16]_i_7__0_n_0 ),
        .I3(\Q[16]_i_8__0_n_0 ),
        .I4(\Q[26]_i_9_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[16]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[16]_i_5__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[13]),
        .I2(STALL_EN),
        .I3(IF_PC2[13]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[13] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[16]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[16]_i_6 
       (.I0(\Q[16]_i_15__0_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[16]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[16]_i_11_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [12]));
  LUT5 #(
    .INIT(32'h02F20EFE)) 
    \Q[16]_i_6__0 
       (.I0(\Q[16]_i_11__0_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [19]),
        .I3(\custom_alu/fp32_add/sel0 [12]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[16]_i_6__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[16]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [16]),
        .O(\Q[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF3FF333F737F737)) 
    \Q[16]_i_7__0 
       (.I0(\Q[26]_i_17_n_0 ),
        .I1(\Q[31]_i_12__0_n_0 ),
        .I2(\Q[17]_i_10__0_n_0 ),
        .I3(\Q[17]_i_15_n_0 ),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[16]_i_7__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[16]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [15]),
        .O(\Q[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEFEEFEFEFFFE)) 
    \Q[16]_i_8__0 
       (.I0(\Q[69]_i_20_n_0 ),
        .I1(\Q[27]_i_13_n_0 ),
        .I2(\Q[28]_i_11_n_0 ),
        .I3(\Q[69]_i_16_n_0 ),
        .I4(\Q[35]_i_28_n_0 ),
        .I5(\Q[35]_i_29_n_0 ),
        .O(\Q[16]_i_8__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[16]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [14]),
        .O(\Q[16]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[16]_i_9__0 
       (.I0(exponent_carry_i_11_n_7),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[16]_i_13_n_4 ),
        .O(\Q[16]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \Q[170]_i_1 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(EX_BR_TAKEN),
        .O(DECODED_INSTRUCTION[0]));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \Q[170]_rep__0_i_1 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(EX_BR_TAKEN),
        .O(\Q[170]_rep__0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \Q[170]_rep__1_i_1 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(EX_BR_TAKEN),
        .O(\Q[170]_rep__1_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \Q[170]_rep__2_i_1 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(EX_BR_TAKEN),
        .O(\Q[170]_rep__2_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \Q[170]_rep__3_i_1 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(EX_BR_TAKEN),
        .O(\Q[170]_rep__3_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \Q[170]_rep_i_1 
       (.I0(I_MEM_DOUT_IBUF[4]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .I5(EX_BR_TAKEN),
        .O(\Q[170]_rep_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFAEAAAE)) 
    \Q[171]_i_1 
       (.I0(\Q[171]_i_2_n_0 ),
        .I1(DECODED_INSTRUCTION[16]),
        .I2(\Q[171]_i_4_n_0 ),
        .I3(\Q[171]_i_5_n_0 ),
        .I4(DECODED_INSTRUCTION[17]),
        .I5(STALL_EN),
        .O(ID_EX_D[171]));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_100 
       (.I0(\Q[47]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[0]),
        .I2(\Q[48]_i_1_n_0 ),
        .I3(ID_RD2_FORWARDED[1]),
        .O(\Q[171]_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[171]_i_101 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[11]),
        .I2(CRF_RD1_IBUF[11]),
        .I3(RF_RD1_IBUF[11]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[171]_i_101_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[171]_i_102 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[9]),
        .I2(CRF_RD1_IBUF[9]),
        .I3(RF_RD1_IBUF[9]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[171]_i_102_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_13 
       (.I0(\Q[78]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[31]),
        .I2(ID_RD2_FORWARDED[30]),
        .I3(\Q[77]_i_1__0_n_0 ),
        .O(\Q[171]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \Q[171]_i_14 
       (.I0(\Q[75]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[28]),
        .I2(\Q[76]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[29]),
        .I4(ID_RD2_FORWARDED[27]),
        .I5(\Q[74]_i_1__0_n_0 ),
        .O(\Q[171]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \Q[171]_i_15 
       (.I0(\Q[73]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[26]),
        .I2(\Q[71]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[24]),
        .I4(\Q[72]_i_1__0_n_0 ),
        .I5(ID_RD2_FORWARDED[25]),
        .O(\Q[171]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[171]_i_17 
       (.I0(ID_RD2_FORWARDED[30]),
        .I1(\Q[77]_i_1__0_n_0 ),
        .O(\Q[171]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_18 
       (.I0(\Q[76]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[29]),
        .I2(ID_RD2_FORWARDED[28]),
        .I3(\Q[75]_i_1__0_n_0 ),
        .O(\Q[171]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_19 
       (.I0(\Q[74]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[27]),
        .I2(ID_RD2_FORWARDED[26]),
        .I3(\Q[73]_i_1__0_n_0 ),
        .O(\Q[171]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEEEEFEEEEEE)) 
    \Q[171]_i_2 
       (.I0(\Q[171]_i_7_n_0 ),
        .I1(ID_JAL_AFTER_LU),
        .I2(\branch_comp/EQ ),
        .I3(\Q[171]_i_9_n_0 ),
        .I4(\Q[90]_i_4_n_0 ),
        .I5(\Q[123]_i_5_n_0 ),
        .O(\Q[171]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_20 
       (.I0(\Q[72]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[25]),
        .I2(ID_RD2_FORWARDED[24]),
        .I3(\Q[71]_i_1__0_n_0 ),
        .O(\Q[171]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \Q[171]_i_21 
       (.I0(ID_RD2_FORWARDED[30]),
        .I1(\Q[77]_i_1__0_n_0 ),
        .O(\Q[171]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_22 
       (.I0(ID_RD2_FORWARDED[29]),
        .I1(\Q[76]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[28]),
        .I3(\Q[75]_i_1__0_n_0 ),
        .O(\Q[171]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_23 
       (.I0(\Q[73]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[26]),
        .I2(ID_RD2_FORWARDED[27]),
        .I3(\Q[74]_i_1__0_n_0 ),
        .O(\Q[171]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_24 
       (.I0(\Q[71]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[24]),
        .I2(\Q[72]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[25]),
        .O(\Q[171]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h2F02)) 
    \Q[171]_i_26 
       (.I0(ID_RD2_FORWARDED[30]),
        .I1(\Q[77]_i_1__0_n_0 ),
        .I2(\Q[78]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[31]),
        .O(\Q[171]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_27 
       (.I0(\Q[76]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[29]),
        .I2(ID_RD2_FORWARDED[28]),
        .I3(\Q[75]_i_1__0_n_0 ),
        .O(\Q[171]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_28 
       (.I0(\Q[74]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[27]),
        .I2(ID_RD2_FORWARDED[26]),
        .I3(\Q[73]_i_1__0_n_0 ),
        .O(\Q[171]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_29 
       (.I0(\Q[72]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[25]),
        .I2(ID_RD2_FORWARDED[24]),
        .I3(\Q[71]_i_1__0_n_0 ),
        .O(\Q[171]_i_29_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    \Q[171]_i_3 
       (.I0(I_MEM_DOUT_IBUF[13]),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .I3(\Q[90]_i_4_n_0 ),
        .O(DECODED_INSTRUCTION[16]));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_30 
       (.I0(\Q[78]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[31]),
        .I2(ID_RD2_FORWARDED[30]),
        .I3(\Q[77]_i_1__0_n_0 ),
        .O(\Q[171]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_31 
       (.I0(ID_RD2_FORWARDED[29]),
        .I1(\Q[76]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[28]),
        .I3(\Q[75]_i_1__0_n_0 ),
        .O(\Q[171]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_32 
       (.I0(\Q[73]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[26]),
        .I2(ID_RD2_FORWARDED[27]),
        .I3(\Q[74]_i_1__0_n_0 ),
        .O(\Q[171]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_33 
       (.I0(\Q[71]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[24]),
        .I2(\Q[72]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[25]),
        .O(\Q[171]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \Q[171]_i_35 
       (.I0(ID_RD2_FORWARDED[23]),
        .I1(\Q[70]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[22]),
        .I3(\Q[69]_i_1__0_n_0 ),
        .I4(ID_RD2_FORWARDED[21]),
        .I5(\Q[68]_i_1__0_n_0 ),
        .O(\Q[171]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \Q[171]_i_36 
       (.I0(ID_RD2_FORWARDED[20]),
        .I1(\Q[67]_i_1__0_n_0 ),
        .I2(\Q[65]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[18]),
        .I4(\Q[66]_i_1__0_n_0 ),
        .I5(ID_RD2_FORWARDED[19]),
        .O(\Q[171]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h00009009)) 
    \Q[171]_i_37 
       (.I0(\Q[63]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[16]),
        .I2(\Q[64]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[17]),
        .I4(\Q[171]_i_61_n_0 ),
        .O(\Q[171]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h41000041)) 
    \Q[171]_i_38 
       (.I0(\Q[171]_i_62_n_0 ),
        .I1(\Q[59]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[12]),
        .I3(\Q[60]_i_1__0_n_0 ),
        .I4(ID_RD2_FORWARDED[13]),
        .O(\Q[171]_i_38_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \Q[171]_i_4 
       (.I0(\Q[90]_i_4_n_0 ),
        .I1(I_MEM_DOUT_IBUF[14]),
        .I2(I_MEM_DOUT_IBUF[13]),
        .O(\Q[171]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hD4)) 
    \Q[171]_i_40 
       (.I0(\Q[70]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[23]),
        .I2(\Q[171]_i_72_n_0 ),
        .O(\Q[171]_i_40_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_41 
       (.I0(\Q[68]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[21]),
        .I2(ID_RD2_FORWARDED[20]),
        .I3(\Q[67]_i_1__0_n_0 ),
        .O(\Q[171]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_42 
       (.I0(\Q[66]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[19]),
        .I2(ID_RD2_FORWARDED[18]),
        .I3(\Q[65]_i_1__0_n_0 ),
        .O(\Q[171]_i_42_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_43 
       (.I0(\Q[64]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[17]),
        .I2(ID_RD2_FORWARDED[16]),
        .I3(\Q[63]_i_1_n_0 ),
        .O(\Q[171]_i_43_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_44 
       (.I0(ID_RD2_FORWARDED[23]),
        .I1(\Q[70]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[22]),
        .I3(\Q[69]_i_1__0_n_0 ),
        .O(\Q[171]_i_44_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_45 
       (.I0(ID_RD2_FORWARDED[20]),
        .I1(\Q[67]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[21]),
        .I3(\Q[68]_i_1__0_n_0 ),
        .O(\Q[171]_i_45_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_46 
       (.I0(\Q[65]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[18]),
        .I2(\Q[66]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[19]),
        .O(\Q[171]_i_46_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_47 
       (.I0(ID_RD2_FORWARDED[17]),
        .I1(\Q[64]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[16]),
        .I3(\Q[63]_i_1_n_0 ),
        .O(\Q[171]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'hD4)) 
    \Q[171]_i_49 
       (.I0(\Q[70]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[23]),
        .I2(\Q[171]_i_72_n_0 ),
        .O(\Q[171]_i_49_n_0 ));
  LUT3 #(
    .INIT(8'hB2)) 
    \Q[171]_i_5 
       (.I0(\Q[78]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[31]),
        .I2(\branch_comp/LT20_in ),
        .O(\Q[171]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_50 
       (.I0(\Q[68]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[21]),
        .I2(ID_RD2_FORWARDED[20]),
        .I3(\Q[67]_i_1__0_n_0 ),
        .O(\Q[171]_i_50_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_51 
       (.I0(\Q[66]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[19]),
        .I2(ID_RD2_FORWARDED[18]),
        .I3(\Q[65]_i_1__0_n_0 ),
        .O(\Q[171]_i_51_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_52 
       (.I0(\Q[64]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[17]),
        .I2(ID_RD2_FORWARDED[16]),
        .I3(\Q[63]_i_1_n_0 ),
        .O(\Q[171]_i_52_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_53 
       (.I0(ID_RD2_FORWARDED[23]),
        .I1(\Q[70]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[22]),
        .I3(\Q[69]_i_1__0_n_0 ),
        .O(\Q[171]_i_53_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_54 
       (.I0(ID_RD2_FORWARDED[20]),
        .I1(\Q[67]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[21]),
        .I3(\Q[68]_i_1__0_n_0 ),
        .O(\Q[171]_i_54_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_55 
       (.I0(\Q[65]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[18]),
        .I2(\Q[66]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[19]),
        .O(\Q[171]_i_55_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_56 
       (.I0(ID_RD2_FORWARDED[17]),
        .I1(\Q[64]_i_1__0_n_0 ),
        .I2(ID_RD2_FORWARDED[16]),
        .I3(\Q[63]_i_1_n_0 ),
        .O(\Q[171]_i_56_n_0 ));
  LUT4 #(
    .INIT(16'h0009)) 
    \Q[171]_i_57 
       (.I0(\Q[57]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[10]),
        .I2(\Q[171]_i_81_n_0 ),
        .I3(\Q[171]_i_82_n_0 ),
        .O(\Q[171]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \Q[171]_i_58 
       (.I0(ID_RD2_FORWARDED[8]),
        .I1(\Q[55]_i_1__0_n_0 ),
        .I2(\Q[53]_i_1_n_0 ),
        .I3(ID_RD2_FORWARDED[6]),
        .I4(\Q[54]_i_1_n_0 ),
        .I5(ID_RD2_FORWARDED[7]),
        .O(\Q[171]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \Q[171]_i_59 
       (.I0(\Q[51]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[4]),
        .I2(\Q[52]_i_1_n_0 ),
        .I3(ID_RD2_FORWARDED[5]),
        .I4(ID_RD2_FORWARDED[3]),
        .I5(\Q[50]_i_1_n_0 ),
        .O(\Q[171]_i_59_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \Q[171]_i_6 
       (.I0(I_MEM_DOUT_IBUF[13]),
        .I1(I_MEM_DOUT_IBUF[14]),
        .I2(I_MEM_DOUT_IBUF[12]),
        .I3(\Q[90]_i_4_n_0 ),
        .O(DECODED_INSTRUCTION[17]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \Q[171]_i_60 
       (.I0(ID_RD2_FORWARDED[2]),
        .I1(\Q[49]_i_1_n_0 ),
        .I2(\Q[47]_i_1_n_0 ),
        .I3(ID_RD2_FORWARDED[0]),
        .I4(\Q[48]_i_1_n_0 ),
        .I5(ID_RD2_FORWARDED[1]),
        .O(\Q[171]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h00000777FFFFF888)) 
    \Q[171]_i_61 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[15]),
        .I2(data0[15]),
        .I3(\Q[78]_i_3_n_0 ),
        .I4(\Q[171]_i_83_n_0 ),
        .I5(ID_RD2_FORWARDED[15]),
        .O(\Q[171]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h00000777FFFFF888)) 
    \Q[171]_i_62 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[14]),
        .I2(data0[14]),
        .I3(\Q[78]_i_3_n_0 ),
        .I4(\Q[171]_i_84_n_0 ),
        .I5(ID_RD2_FORWARDED[14]),
        .O(\Q[171]_i_62_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_64 
       (.I0(\Q[62]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[15]),
        .I2(ID_RD2_FORWARDED[14]),
        .I3(\Q[61]_i_1__0_n_0 ),
        .O(\Q[171]_i_64_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_65 
       (.I0(\Q[60]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[13]),
        .I2(ID_RD2_FORWARDED[12]),
        .I3(\Q[59]_i_1__0_n_0 ),
        .O(\Q[171]_i_65_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_66 
       (.I0(\Q[58]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[11]),
        .I2(ID_RD2_FORWARDED[10]),
        .I3(\Q[57]_i_1__0_n_0 ),
        .O(\Q[171]_i_66_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_67 
       (.I0(\Q[56]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[9]),
        .I2(ID_RD2_FORWARDED[8]),
        .I3(\Q[55]_i_1__0_n_0 ),
        .O(\Q[171]_i_67_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \Q[171]_i_68 
       (.I0(\Q[171]_i_62_n_0 ),
        .I1(\Q[171]_i_61_n_0 ),
        .O(\Q[171]_i_68_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_69 
       (.I0(\Q[59]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[12]),
        .I2(\Q[60]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[13]),
        .O(\Q[171]_i_69_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT5 #(
    .INIT(32'h60000000)) 
    \Q[171]_i_7 
       (.I0(\Q_reg[171]_i_11_n_0 ),
        .I1(I_MEM_DOUT_IBUF[12]),
        .I2(I_MEM_DOUT_IBUF[13]),
        .I3(I_MEM_DOUT_IBUF[14]),
        .I4(\Q[90]_i_4_n_0 ),
        .O(\Q[171]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h41)) 
    \Q[171]_i_70 
       (.I0(\Q[171]_i_81_n_0 ),
        .I1(ID_RD2_FORWARDED[10]),
        .I2(\Q[57]_i_1__0_n_0 ),
        .O(\Q[171]_i_70_n_0 ));
  LUT3 #(
    .INIT(8'h09)) 
    \Q[171]_i_71 
       (.I0(ID_RD2_FORWARDED[8]),
        .I1(\Q[55]_i_1__0_n_0 ),
        .I2(\Q[171]_i_82_n_0 ),
        .O(\Q[171]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFF888)) 
    \Q[171]_i_72 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(data1[22]),
        .I2(data0[22]),
        .I3(\Q[46]_i_3_n_0 ),
        .I4(\Q[37]_i_2_n_0 ),
        .I5(\Q[69]_i_1__0_n_0 ),
        .O(\Q[171]_i_72_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_74 
       (.I0(\Q[60]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[13]),
        .I2(ID_RD2_FORWARDED[12]),
        .I3(\Q[59]_i_1__0_n_0 ),
        .O(\Q[171]_i_74_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_75 
       (.I0(\Q[58]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[11]),
        .I2(ID_RD2_FORWARDED[10]),
        .I3(\Q[57]_i_1__0_n_0 ),
        .O(\Q[171]_i_75_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_76 
       (.I0(\Q[56]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[9]),
        .I2(ID_RD2_FORWARDED[8]),
        .I3(\Q[55]_i_1__0_n_0 ),
        .O(\Q[171]_i_76_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \Q[171]_i_77 
       (.I0(\Q[171]_i_62_n_0 ),
        .I1(\Q[171]_i_61_n_0 ),
        .O(\Q[171]_i_77_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_78 
       (.I0(\Q[59]_i_1__0_n_0 ),
        .I1(ID_RD2_FORWARDED[12]),
        .I2(\Q[60]_i_1__0_n_0 ),
        .I3(ID_RD2_FORWARDED[13]),
        .O(\Q[171]_i_78_n_0 ));
  LUT3 #(
    .INIT(8'h41)) 
    \Q[171]_i_79 
       (.I0(\Q[171]_i_81_n_0 ),
        .I1(ID_RD2_FORWARDED[10]),
        .I2(\Q[57]_i_1__0_n_0 ),
        .O(\Q[171]_i_79_n_0 ));
  LUT3 #(
    .INIT(8'h09)) 
    \Q[171]_i_80 
       (.I0(ID_RD2_FORWARDED[8]),
        .I1(\Q[55]_i_1__0_n_0 ),
        .I2(\Q[171]_i_82_n_0 ),
        .O(\Q[171]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h00000777FFFFF888)) 
    \Q[171]_i_81 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[11]),
        .I2(data0[11]),
        .I3(\Q[78]_i_3_n_0 ),
        .I4(\Q[171]_i_101_n_0 ),
        .I5(ID_RD2_FORWARDED[11]),
        .O(\Q[171]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h00000777FFFFF888)) 
    \Q[171]_i_82 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[9]),
        .I2(data0[9]),
        .I3(\Q[78]_i_3_n_0 ),
        .I4(\Q[171]_i_102_n_0 ),
        .I5(ID_RD2_FORWARDED[9]),
        .O(\Q[171]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[171]_i_83 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[15]),
        .I2(CRF_RD1_IBUF[15]),
        .I3(RF_RD1_IBUF[15]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[171]_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[171]_i_84 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[14]),
        .I2(CRF_RD1_IBUF[14]),
        .I3(RF_RD1_IBUF[14]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[171]_i_84_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_85 
       (.I0(\Q[54]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[7]),
        .I2(ID_RD2_FORWARDED[6]),
        .I3(\Q[53]_i_1_n_0 ),
        .O(\Q[171]_i_85_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_86 
       (.I0(\Q[52]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[5]),
        .I2(ID_RD2_FORWARDED[4]),
        .I3(\Q[51]_i_1_n_0 ),
        .O(\Q[171]_i_86_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_87 
       (.I0(\Q[50]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[3]),
        .I2(ID_RD2_FORWARDED[2]),
        .I3(\Q[49]_i_1_n_0 ),
        .O(\Q[171]_i_87_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_88 
       (.I0(\Q[48]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[1]),
        .I2(ID_RD2_FORWARDED[0]),
        .I3(\Q[47]_i_1_n_0 ),
        .O(\Q[171]_i_88_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_89 
       (.I0(\Q[53]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[6]),
        .I2(\Q[54]_i_1_n_0 ),
        .I3(ID_RD2_FORWARDED[7]),
        .O(\Q[171]_i_89_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \Q[171]_i_9 
       (.I0(I_MEM_DOUT_IBUF[12]),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[14]),
        .O(\Q[171]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_90 
       (.I0(ID_RD2_FORWARDED[5]),
        .I1(\Q[52]_i_1_n_0 ),
        .I2(ID_RD2_FORWARDED[4]),
        .I3(\Q[51]_i_1_n_0 ),
        .O(\Q[171]_i_90_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_91 
       (.I0(ID_RD2_FORWARDED[2]),
        .I1(\Q[49]_i_1_n_0 ),
        .I2(ID_RD2_FORWARDED[3]),
        .I3(\Q[50]_i_1_n_0 ),
        .O(\Q[171]_i_91_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_92 
       (.I0(\Q[47]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[0]),
        .I2(\Q[48]_i_1_n_0 ),
        .I3(ID_RD2_FORWARDED[1]),
        .O(\Q[171]_i_92_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_93 
       (.I0(\Q[54]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[7]),
        .I2(ID_RD2_FORWARDED[6]),
        .I3(\Q[53]_i_1_n_0 ),
        .O(\Q[171]_i_93_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_94 
       (.I0(\Q[52]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[5]),
        .I2(ID_RD2_FORWARDED[4]),
        .I3(\Q[51]_i_1_n_0 ),
        .O(\Q[171]_i_94_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_95 
       (.I0(\Q[50]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[3]),
        .I2(ID_RD2_FORWARDED[2]),
        .I3(\Q[49]_i_1_n_0 ),
        .O(\Q[171]_i_95_n_0 ));
  LUT4 #(
    .INIT(16'h44D4)) 
    \Q[171]_i_96 
       (.I0(\Q[48]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[1]),
        .I2(ID_RD2_FORWARDED[0]),
        .I3(\Q[47]_i_1_n_0 ),
        .O(\Q[171]_i_96_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_97 
       (.I0(\Q[53]_i_1_n_0 ),
        .I1(ID_RD2_FORWARDED[6]),
        .I2(\Q[54]_i_1_n_0 ),
        .I3(ID_RD2_FORWARDED[7]),
        .O(\Q[171]_i_97_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_98 
       (.I0(ID_RD2_FORWARDED[5]),
        .I1(\Q[52]_i_1_n_0 ),
        .I2(ID_RD2_FORWARDED[4]),
        .I3(\Q[51]_i_1_n_0 ),
        .O(\Q[171]_i_98_n_0 ));
  LUT4 #(
    .INIT(16'h9009)) 
    \Q[171]_i_99 
       (.I0(ID_RD2_FORWARDED[2]),
        .I1(\Q[49]_i_1_n_0 ),
        .I2(ID_RD2_FORWARDED[3]),
        .I3(\Q[50]_i_1_n_0 ),
        .O(\Q[171]_i_99_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[17]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [17]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [16]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [17]));
  LUT6 #(
    .INIT(64'h1111100000001000)) 
    \Q[17]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [11]),
        .I2(\custom_alu/fp32_add/sel0 [8]),
        .I3(\custom_alu/fp32_add/sel0 [2]),
        .I4(\custom_alu/fp32_add/sel0 [9]),
        .I5(\custom_alu/fp32_add/sel0 [3]),
        .O(\Q[17]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[17]_i_10__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [16]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[142]),
        .I5(EX_RF_RD1[16]),
        .O(\Q[17]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAACC00AAAACC0F)) 
    \Q[17]_i_11 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [4]),
        .I2(\Q[17]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [10]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .I5(\Q[17]_i_13_n_0 ),
        .O(\Q[17]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[17]_i_11__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [14]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[140]),
        .I5(EX_RF_RD1[14]),
        .O(\Q[17]_i_11__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT4 #(
    .INIT(16'h4777)) 
    \Q[17]_i_12 
       (.I0(\custom_alu/fp32_add/sel0 [1]),
        .I1(\custom_alu/fp32_add/sel0 [7]),
        .I2(\custom_alu/fp32_add/sel0 [0]),
        .I3(\custom_alu/fp32_add/sel0 [6]),
        .O(\Q[17]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \Q[17]_i_12__0 
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[152]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [26]),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[17]_i_12__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \Q[17]_i_13 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [9]),
        .O(\Q[17]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBABBAAAABABB)) 
    \Q[17]_i_13__0 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[17]_i_19_n_0 ),
        .I2(\Q[21]_i_10__0_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[67]_i_12_n_0 ),
        .I5(\Q[17]_i_20_n_0 ),
        .O(\Q[17]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[17]_i_14 
       (.I0(\custom_alu/int2fp/INT_VAL0 [15]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[141]),
        .I5(EX_RF_RD1[15]),
        .O(\Q[17]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[17]_i_15 
       (.I0(\custom_alu/int2fp/INT_VAL0 [4]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[130]),
        .I5(EX_RF_RD1[4]),
        .O(\Q[17]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \Q[17]_i_16 
       (.I0(\Q[28]_i_18_n_0 ),
        .I1(\Q[35]_i_32_n_0 ),
        .I2(\Q[17]_i_21_n_0 ),
        .I3(\Q[17]_i_11__0_n_0 ),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[17]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0004FF0400F4FFF4)) 
    \Q[17]_i_17 
       (.I0(\Q[35]_i_28_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[35]_i_26_n_0 ),
        .I5(\Q[35]_i_29_n_0 ),
        .O(\Q[17]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00000777)) 
    \Q[17]_i_18 
       (.I0(\Q[28]_i_7_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[28]_i_11_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .O(\Q[17]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB800B800B800)) 
    \Q[17]_i_19 
       (.I0(\custom_alu/int2fp/INT_VAL0 [10]),
        .I1(PSUM3__0_carry__0_i_10__2_n_0),
        .I2(ALU_DIN1[10]),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[31]_i_11__0_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[17]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[17]_i_1__0 
       (.I0(\Q[17]_i_2_n_0 ),
        .I1(\Q[17]_i_3_n_0 ),
        .I2(\Q[17]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[18] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [17]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[17]_i_1__1 
       (.I0(\Q[17]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[2]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[2]),
        .I5(\Q[17]_i_3__1_n_0 ),
        .O(ID_RD2_FORWARDED[2]));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \Q[17]_i_1__2 
       (.I0(\Q[17]_i_2__0_n_0 ),
        .I1(\Q[17]_i_3__0_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\Q[17]_i_4__0_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[12]),
        .O(data0[12]));
  LUT6 #(
    .INIT(64'hFFFFF8FF0000F800)) 
    \Q[17]_i_1__3 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(\Q[17]_i_2__2_n_0 ),
        .I3(EX_MEM_Q[39]),
        .I4(EX_MEM_Q[37]),
        .I5(EX_MEM_Q[17]),
        .O(data1[12]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[17]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [17]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [17]),
        .O(\Q[17]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h30353F35)) 
    \Q[17]_i_20 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[28]_i_18_n_0 ),
        .I2(\Q[29]_i_10_n_0 ),
        .I3(\Q[28]_i_20_n_0 ),
        .I4(\Q[35]_i_20_n_0 ),
        .O(\Q[17]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8888888B888)) 
    \Q[17]_i_21 
       (.I0(\Q[47]_i_9_n_0 ),
        .I1(\Q[35]_i_20_n_0 ),
        .I2(\Q[35]_i_19_n_0 ),
        .I3(EX_RF_RD1[0]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I5(ID_EX_Q[126]),
        .O(\Q[17]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h2222222220200020)) 
    \Q[17]_i_2__0 
       (.I0(\Q[17]_i_5__0_n_0 ),
        .I1(\Q[17]_i_6__0_n_0 ),
        .I2(\Q[26]_i_7_n_0 ),
        .I3(\Q[17]_i_7__0_n_0 ),
        .I4(\Q[17]_i_8__0_n_0 ),
        .I5(\Q[17]_i_9__0_n_0 ),
        .O(\Q[17]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[17]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[2]),
        .I2(CRF_RD2_IBUF[2]),
        .I3(RF_RD2_IBUF[2]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[17]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AA8080000A808)) 
    \Q[17]_i_2__2 
       (.I0(\Q[11]_i_5__1_n_0 ),
        .I1(D_MEM_DOUT_IBUF[12]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I3(D_MEM_DOUT_IBUF[28]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[20]),
        .O(\Q[17]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFFDCDFCCCFDCD)) 
    \Q[17]_i_3 
       (.I0(\Q[17]_i_5_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [21]),
        .I3(\custom_alu/fp32_add/sel0 [15]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [14]),
        .O(\Q[17]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[17]_i_3__0 
       (.I0(\custom_alu/fp32_mult/product_mantissa [12]),
        .I1(\Q[65]_i_5_n_0 ),
        .O(\Q[17]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[17]_i_3__1 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(data1[2]),
        .O(\Q[17]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT4 #(
    .INIT(16'hF4FF)) 
    \Q[17]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [16]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [23]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB8B8888BB8B)) 
    \Q[17]_i_4__0 
       (.I0(\custom_alu/MULT [12]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(EX_CUSTOM_ALU_SEL[29]),
        .I3(\custom_alu/Q [12]),
        .I4(EX_CUSTOM_ALU_SEL[30]),
        .I5(\custom_alu/MULT [44]),
        .O(\Q[17]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT5 #(
    .INIT(32'h02F20EFE)) 
    \Q[17]_i_5 
       (.I0(\Q[17]_i_6_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [19]),
        .I3(\custom_alu/fp32_add/sel0 [13]),
        .I4(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[17]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEFEAFFFF)) 
    \Q[17]_i_5__0 
       (.I0(INT0_carry__1_i_5_n_0),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[17]_i_5__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[17]_i_6 
       (.I0(\custom_alu/fp32_add/sel0 [11]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [10]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\Q[17]_i_7_n_0 ),
        .O(\Q[17]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[17]_i_6__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [12]),
        .O(\Q[17]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h7474747774747444)) 
    \Q[17]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [9]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\Q[17]_i_8_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [13]),
        .I4(\custom_alu/fp32_add/sel0 [14]),
        .I5(\Q[17]_i_9_n_0 ),
        .O(\Q[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5555003F55550000)) 
    \Q[17]_i_7__0 
       (.I0(\Q[17]_i_10__0_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[17]_i_12__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[17]_i_13__0_n_0 ),
        .O(\Q[17]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \Q[17]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [14]),
        .I2(\custom_alu/fp32_add/sel0 [7]),
        .O(\Q[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FFD5)) 
    \Q[17]_i_8__0 
       (.I0(\Q[22]_i_7__0_n_0 ),
        .I1(\Q[17]_i_14_n_0 ),
        .I2(\Q[17]_i_15_n_0 ),
        .I3(\Q[17]_i_16_n_0 ),
        .I4(\Q[17]_i_17_n_0 ),
        .I5(\Q[27]_i_13_n_0 ),
        .O(\Q[17]_i_8__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT4 #(
    .INIT(16'h4447)) 
    \Q[17]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .I2(\Q[17]_i_10_n_0 ),
        .I3(\Q[17]_i_11_n_0 ),
        .O(\Q[17]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF4540FFFFFFFF)) 
    \Q[17]_i_9__0 
       (.I0(\Q[17]_i_18_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[28]_i_6_n_0 ),
        .I3(\Q[26]_i_15__0_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[17]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[18]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [18]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [17]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [18]));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT5 #(
    .INIT(32'hFFFFF808)) 
    \Q[18]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [5]),
        .I2(\custom_alu/fp32_add/sel0 [11]),
        .I3(\custom_alu/fp32_add/sel0 [6]),
        .I4(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[18]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h0000CAC0)) 
    \Q[18]_i_10__0 
       (.I0(\Q[29]_i_18__0_n_0 ),
        .I1(\Q[17]_i_15_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[28]_i_18_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .O(\Q[18]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'hFF00B8B800000000)) 
    \Q[18]_i_11 
       (.I0(\custom_alu/fp32_add/sel0 [3]),
        .I1(\custom_alu/fp32_add/sel0 [8]),
        .I2(\Q[18]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [4]),
        .I4(\custom_alu/fp32_add/sel0 [9]),
        .I5(exp_sub_carry__0_i_6_n_0),
        .O(\Q[18]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \Q[18]_i_11__0 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[17]_i_14_n_0 ),
        .I4(\Q[35]_i_28_n_0 ),
        .O(\Q[18]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[18]_i_12 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [7]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [6]),
        .I4(\custom_alu/fp32_add/sel0 [5]),
        .I5(\custom_alu/fp32_add/sel0 [0]),
        .O(\Q[18]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF088)) 
    \Q[18]_i_12__0 
       (.I0(\Q[35]_i_21_n_0 ),
        .I1(ALU_DIN1[0]),
        .I2(\Q[47]_i_9_n_0 ),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[35]_i_20_n_0 ),
        .O(\Q[18]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0FFFFFFF1FFF1)) 
    \Q[18]_i_13 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[35]_i_21_n_0 ),
        .I2(\Q[17]_i_14_n_0 ),
        .I3(\Q[35]_i_24_n_0 ),
        .I4(\Q[35]_i_32_n_0 ),
        .I5(\Q[35]_i_20_n_0 ),
        .O(\Q[18]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00040F04F0F4FFF4)) 
    \Q[18]_i_14 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[28]_i_11_n_0 ),
        .I3(\Q[69]_i_16_n_0 ),
        .I4(\Q[35]_i_26_n_0 ),
        .I5(\Q[35]_i_27_n_0 ),
        .O(\Q[18]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8B8B88B888888)) 
    \Q[18]_i_15 
       (.I0(\Q[17]_i_11__0_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[35]_i_20_n_0 ),
        .I4(\Q[31]_i_13__0_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[18]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000F77FFFF0F77)) 
    \Q[18]_i_16 
       (.I0(\Q[35]_i_22_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[35]_i_21_n_0 ),
        .I3(\Q[31]_i_11__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[35]_i_19_n_0 ),
        .O(\Q[18]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \Q[18]_i_17 
       (.I0(\Q[17]_i_14_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[17]_i_10__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[18]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[18]_i_1__0 
       (.I0(\Q[18]_i_2_n_0 ),
        .I1(\Q[18]_i_3_n_0 ),
        .I2(\Q[18]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[19] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [18]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[18]_i_1__1 
       (.I0(\Q[18]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[3]),
        .I3(data1[3]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[3]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[18]_i_1__2 
       (.I0(\Q[18]_i_2__0_n_0 ),
        .I1(\Q[18]_i_3__0_n_0 ),
        .I2(\Q[18]_i_4__0_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[13]),
        .O(data0[13]));
  LUT6 #(
    .INIT(64'hFFFFF8FF0000F800)) 
    \Q[18]_i_1__3 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(\Q[18]_i_2__2_n_0 ),
        .I3(EX_MEM_Q[39]),
        .I4(EX_MEM_Q[37]),
        .I5(EX_MEM_Q[18]),
        .O(data1[13]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[18]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [18]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [18]),
        .O(\Q[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[18]_i_2__0 
       (.I0(\custom_alu/MULT [13]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [45]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [13]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[18]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[18]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[3]),
        .I2(CRF_RD2_IBUF[3]),
        .I3(RF_RD2_IBUF[3]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[18]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AA8080000A808)) 
    \Q[18]_i_2__2 
       (.I0(\Q[11]_i_5__1_n_0 ),
        .I1(D_MEM_DOUT_IBUF[13]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I3(D_MEM_DOUT_IBUF[29]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[21]),
        .O(\Q[18]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFFCDDFCCCFCDD)) 
    \Q[18]_i_3 
       (.I0(\Q[18]_i_5_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [16]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [15]),
        .O(\Q[18]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \Q[18]_i_3__0 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [13]),
        .O(\Q[18]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT4 #(
    .INIT(16'hBBFB)) 
    \Q[18]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [23]),
        .I1(\custom_alu/fp32_add/sel0 [24]),
        .I2(\custom_alu/fp32_add/sel0 [22]),
        .I3(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3233023332000200)) 
    \Q[18]_i_4__0 
       (.I0(INT0_carry__2_i_9_n_0),
        .I1(EX_CUSTOM_ALU_SEL[28]),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(EX_CUSTOM_ALU_SEL[27]),
        .I4(\custom_alu/fp2int/INT0 [13]),
        .I5(\Q[18]_i_5__0_n_0 ),
        .O(\Q[18]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT5 #(
    .INIT(32'h02F20EFE)) 
    \Q[18]_i_5 
       (.I0(\Q[18]_i_6_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [19]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\custom_alu/fp32_add/sel0 [13]),
        .O(\Q[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAAA88888888)) 
    \Q[18]_i_5__0 
       (.I0(EX_CUSTOM_ALU_SEL[26]),
        .I1(\Q[18]_i_6__0_n_0 ),
        .I2(\Q[18]_i_7__0_n_0 ),
        .I3(\Q[18]_i_8__0_n_0 ),
        .I4(\Q[18]_i_9__0_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[18]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h5554FFFF55545554)) 
    \Q[18]_i_6 
       (.I0(\Q[18]_i_7_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [16]),
        .I2(\custom_alu/fp32_add/sel0 [15]),
        .I3(\Q[18]_i_8_n_0 ),
        .I4(\custom_alu/fp32_add/sel0 [12]),
        .I5(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[18]_i_6__0 
       (.I0(\Q[31]_i_11__0_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[31]_i_10__0_n_0 ),
        .I4(\Q[28]_i_11_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[18]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF088)) 
    \Q[18]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [11]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \Q[18]_i_7__0 
       (.I0(EX_RF_RD1[17]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[143]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [17]),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[18]_i_7__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT5 #(
    .INIT(32'h553F5530)) 
    \Q[18]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [9]),
        .I1(\custom_alu/fp32_add/sel0 [8]),
        .I2(\custom_alu/fp32_add/sel0 [13]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\Q[18]_i_9_n_0 ),
        .O(\Q[18]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000EEFE)) 
    \Q[18]_i_8__0 
       (.I0(\Q[18]_i_10__0_n_0 ),
        .I1(\Q[18]_i_11__0_n_0 ),
        .I2(\Q[18]_i_12__0_n_0 ),
        .I3(\Q[18]_i_13_n_0 ),
        .I4(\Q[18]_i_14_n_0 ),
        .I5(\Q[27]_i_13_n_0 ),
        .O(\Q[18]_i_8__0_n_0 ));
  LUT4 #(
    .INIT(16'h444F)) 
    \Q[18]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .I2(\Q[18]_i_10_n_0 ),
        .I3(\Q[18]_i_11_n_0 ),
        .O(\Q[18]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1110)) 
    \Q[18]_i_9__0 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[18]_i_15_n_0 ),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[18]_i_16_n_0 ),
        .I4(\Q[18]_i_17_n_0 ),
        .O(\Q[18]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[19]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [19]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [18]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [19]));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT5 #(
    .INIT(32'hFFFFF808)) 
    \Q[19]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [6]),
        .I2(\custom_alu/fp32_add/sel0 [11]),
        .I3(\custom_alu/fp32_add/sel0 [7]),
        .I4(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[19]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EFEEEFFF)) 
    \Q[19]_i_11 
       (.I0(\custom_alu/fp32_add/sel0 [9]),
        .I1(\custom_alu/fp32_add/sel0 [8]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [7]),
        .I4(\Q[19]_i_12_n_0 ),
        .I5(\Q[19]_i_13_n_0 ),
        .O(\Q[19]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[19]_i_12 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [6]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [5]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [4]),
        .O(\Q[19]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hB888)) 
    \Q[19]_i_13 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [9]),
        .I2(\custom_alu/fp32_add/sel0 [4]),
        .I3(\custom_alu/fp32_add/sel0 [8]),
        .O(\Q[19]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[19]_i_1__0 
       (.I0(\Q[19]_i_2_n_0 ),
        .I1(\Q[19]_i_3_n_0 ),
        .I2(\Q[19]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[20] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [19]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[19]_i_1__1 
       (.I0(\Q[19]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[4]),
        .I3(data1[4]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[4]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[19]_i_1__2 
       (.I0(\Q[19]_i_2__0_n_0 ),
        .I1(\Q[34]_i_5_n_0 ),
        .I2(\Q[19]_i_3__0_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[14]),
        .O(data0[14]));
  LUT6 #(
    .INIT(64'hFFFFF8FF0000F800)) 
    \Q[19]_i_1__3 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(\Q[19]_i_3__1_n_0 ),
        .I3(EX_MEM_Q[39]),
        .I4(EX_MEM_Q[37]),
        .I5(EX_MEM_Q[19]),
        .O(data1[14]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[19]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [19]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [19]),
        .O(\Q[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0B00FFFF0B000B00)) 
    \Q[19]_i_2__0 
       (.I0(\Q[19]_i_4__0_n_0 ),
        .I1(\Q[19]_i_5__0_n_0 ),
        .I2(\Q[29]_i_6__0_n_0 ),
        .I3(\Q[29]_i_7__0_n_0 ),
        .I4(\Q[65]_i_5_n_0 ),
        .I5(\custom_alu/fp32_mult/product_mantissa [14]),
        .O(\Q[19]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[19]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[4]),
        .I2(CRF_RD2_IBUF[4]),
        .I3(RF_RD2_IBUF[4]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[19]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[19]_i_2__2 
       (.I0(D_MEM_DOUT_IBUF[15]),
        .I1(D_MEM_DOUT_IBUF[7]),
        .I2(D_MEM_DOUT_IBUF[31]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[23]),
        .O(\Q[19]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFFCDDFCCCFCDD)) 
    \Q[19]_i_3 
       (.I0(\Q[19]_i_5_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [17]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [16]),
        .O(\Q[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB8B8888BB8B)) 
    \Q[19]_i_3__0 
       (.I0(\custom_alu/MULT [14]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(EX_CUSTOM_ALU_SEL[29]),
        .I3(\custom_alu/Q [14]),
        .I4(EX_CUSTOM_ALU_SEL[30]),
        .I5(\custom_alu/MULT [46]),
        .O(\Q[19]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AA8080000A808)) 
    \Q[19]_i_3__1 
       (.I0(\Q[11]_i_5__1_n_0 ),
        .I1(D_MEM_DOUT_IBUF[14]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I3(D_MEM_DOUT_IBUF[30]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[22]),
        .O(\Q[19]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT4 #(
    .INIT(16'hBBFB)) 
    \Q[19]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [23]),
        .I1(\custom_alu/fp32_add/sel0 [24]),
        .I2(\custom_alu/fp32_add/sel0 [22]),
        .I3(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF4540FFFFFFFF)) 
    \Q[19]_i_4__0 
       (.I0(\Q[19]_i_7__0_n_0 ),
        .I1(\Q[31]_i_14__0_n_0 ),
        .I2(\Q[28]_i_6_n_0 ),
        .I3(\Q[26]_i_15__0_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[19]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFEEFE)) 
    \Q[19]_i_5 
       (.I0(\custom_alu/fp32_add/sel0 [19]),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [17]),
        .I3(\custom_alu/fp32_add/sel0 [13]),
        .I4(\Q[19]_i_6_n_0 ),
        .I5(\Q[19]_i_7_n_0 ),
        .O(\Q[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h70770000FFFFFFFF)) 
    \Q[19]_i_5__0 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(\Q[28]_i_11_n_0 ),
        .I2(\Q[29]_i_11_n_0 ),
        .I3(\Q[29]_i_10__0_n_0 ),
        .I4(\Q[29]_i_9_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[19]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0030023203330232)) 
    \Q[19]_i_6 
       (.I0(\Q[19]_i_8_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [16]),
        .I3(\custom_alu/fp32_add/sel0 [12]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[19]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT4 #(
    .INIT(16'hB888)) 
    \Q[19]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [15]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [14]),
        .I3(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[19]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00000777)) 
    \Q[19]_i_7__0 
       (.I0(\Q[28]_i_7_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .O(\Q[19]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h553F5530)) 
    \Q[19]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [9]),
        .I2(\custom_alu/fp32_add/sel0 [13]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\Q[19]_i_9_n_0 ),
        .O(\Q[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4F4F4F4F44)) 
    \Q[19]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .I2(\Q[19]_i_10_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [10]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .I5(\Q[19]_i_11_n_0 ),
        .O(\Q[19]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[1]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [0]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [1]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [1]));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT4 #(
    .INIT(16'h0454)) 
    \Q[1]_i_1__0 
       (.I0(\Q[31]_i_2__1_n_0 ),
        .I1(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[2] ),
        .I2(\Q[30]_i_2__1_n_0 ),
        .I3(\Q[1]_i_2_n_0 ),
        .O(\custom_alu/FADD_Q [1]));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[1]_i_1__1 
       (.I0(I_MEM_DOUT_IBUF[8]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[8]));
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'h14)) 
    \Q[1]_i_1__2 
       (.I0(STALL_COUNTER_D1),
        .I1(STALL_COUNTER_Q[0]),
        .I2(STALL_COUNTER_Q[1]),
        .O(STALL_COUNTER_D[1]));
  LUT6 #(
    .INIT(64'h303F3F3F55555555)) 
    \Q[1]_i_2 
       (.I0(\custom_alu/fp32_add/data23 [1]),
        .I1(\custom_alu/fp32_add/sel0 [1]),
        .I2(\custom_alu/fp32_add/sel0 [23]),
        .I3(\custom_alu/fp32_add/sel0 [0]),
        .I4(\custom_alu/fp32_add/sel0 [22]),
        .I5(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[1]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[20]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [20]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [19]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [20]));
  LUT5 #(
    .INIT(32'hFFFFF808)) 
    \Q[20]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [7]),
        .I2(\custom_alu/fp32_add/sel0 [11]),
        .I3(\custom_alu/fp32_add/sel0 [8]),
        .I4(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[20]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[20]_i_10__0 
       (.I0(exponent_carry_i_11_n_4),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_11_n_5),
        .O(\Q[20]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h54FF5454FFFFFFFF)) 
    \Q[20]_i_11 
       (.I0(\Q[20]_i_12_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [8]),
        .I2(\Q[20]_i_13_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [6]),
        .I4(\custom_alu/fp32_add/sel0 [9]),
        .I5(exp_sub_carry__0_i_6_n_0),
        .O(\Q[20]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[20]_i_11__0 
       (.I0(exponent_carry_i_11_n_5),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_11_n_6),
        .O(\Q[20]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h0303000023202320)) 
    \Q[20]_i_11__1 
       (.I0(\Q[23]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[20]_i_19_n_0 ),
        .I4(\Q[23]_i_19_n_0 ),
        .I5(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[20]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF001000)) 
    \Q[20]_i_12 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [6]),
        .I2(\custom_alu/fp32_add/sel0 [2]),
        .I3(\custom_alu/fp32_add/sel0 [5]),
        .I4(\custom_alu/fp32_add/sel0 [8]),
        .I5(\custom_alu/fp32_add/sel0 [9]),
        .O(\Q[20]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[20]_i_12__0 
       (.I0(exponent_carry_i_11_n_6),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_11_n_7),
        .O(\Q[20]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h0033000000B800B8)) 
    \Q[20]_i_12__1 
       (.I0(\Q[23]_i_20_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[20]_i_20_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I4(\Q[23]_i_21_n_0 ),
        .I5(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[20]_i_12__1_n_0 ));
  LUT6 #(
    .INIT(64'h0A0AAAAA0A0A8AAA)) 
    \Q[20]_i_13 
       (.I0(\Q[20]_i_14__0_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [5]),
        .I2(\custom_alu/fp32_add/sel0 [4]),
        .I3(\custom_alu/fp32_add/sel0 [1]),
        .I4(\custom_alu/fp32_add/sel0 [7]),
        .I5(\custom_alu/fp32_add/sel0 [6]),
        .O(\Q[20]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000F44FFFF0F44)) 
    \Q[20]_i_13__0 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[35]_i_22_n_0 ),
        .I3(\Q[69]_i_16_n_0 ),
        .I4(\Q[28]_i_11_n_0 ),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[20]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h2320FFFF23200000)) 
    \Q[20]_i_13__1 
       (.I0(\Q[23]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[20]_i_19_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I5(\Q[16]_i_12_n_0 ),
        .O(\Q[20]_i_13__1_n_0 ));
  LUT5 #(
    .INIT(32'h002AAA2A)) 
    \Q[20]_i_14 
       (.I0(\Q[69]_i_20_n_0 ),
        .I1(ALU_DIN1[0]),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[47]_i_9_n_0 ),
        .O(\Q[20]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FFEFFFFFFFFF)) 
    \Q[20]_i_14__0 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [5]),
        .I2(\custom_alu/fp32_add/sel0 [0]),
        .I3(\custom_alu/fp32_add/sel0 [7]),
        .I4(\custom_alu/fp32_add/sel0 [6]),
        .I5(\custom_alu/fp32_add/sel0 [3]),
        .O(\Q[20]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \Q[20]_i_14__1 
       (.I0(\Q[23]_i_20_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[20]_i_20_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I5(\Q[20]_i_21_n_0 ),
        .O(\Q[20]_i_14__1_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[20]_i_15 
       (.I0(ID_EX_Q[98]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[19]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[19]),
        .O(\Q[20]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[20]_i_16 
       (.I0(ID_EX_Q[97]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[18]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[18]),
        .O(\Q[20]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[20]_i_17 
       (.I0(ID_EX_Q[96]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[17]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[17]),
        .O(\Q[20]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[20]_i_18 
       (.I0(ID_EX_Q[95]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[16]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[16]),
        .O(\Q[20]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[20]_i_19 
       (.I0(EX_RF_RD2[19]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[98]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[19]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[20]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[20]_i_1__0 
       (.I0(\Q[20]_i_2_n_0 ),
        .I1(\Q[20]_i_3__0_n_0 ),
        .I2(\Q[20]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[21] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [20]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[20]_i_1__1 
       (.I0(\Q[20]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[5]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[5]),
        .I5(\Q[20]_i_3__2_n_0 ),
        .O(ID_RD2_FORWARDED[5]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[20]_i_1__2 
       (.I0(\Q[20]_i_2__0_n_0 ),
        .I1(\Q[20]_i_3__1_n_0 ),
        .I2(\Q[20]_i_4__1_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[15]),
        .O(data0[15]));
  LUT6 #(
    .INIT(64'hAAAAEEEEAAFAEEEE)) 
    \Q[20]_i_1__3 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[20]),
        .I2(\Q[20]_i_2__2_n_0 ),
        .I3(MEM_LOAD_SEL[2]),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(\Q[20]_i_4__2_n_0 ),
        .O(data1[15]));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[20]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [20]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [20]),
        .O(\Q[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[20]_i_20 
       (.I0(EX_RF_RD2[18]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[97]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[18]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[20]_i_20_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[20]_i_21 
       (.I0(\Q[23]_i_21_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[20]_i_22_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [3]),
        .O(\Q[20]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[20]_i_22 
       (.I0(EX_RF_RD2[16]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[95]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[16]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[20]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[20]_i_2__0 
       (.I0(\custom_alu/MULT [15]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [47]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [15]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[20]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[20]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[5]),
        .I2(CRF_RD2_IBUF[5]),
        .I3(RF_RD2_IBUF[5]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[20]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \Q[20]_i_2__2 
       (.I0(D_MEM_DOUT_IBUF[23]),
        .I1(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I2(D_MEM_DOUT_IBUF[31]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(D_MEM_DOUT_IBUF[15]),
        .O(\Q[20]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[20]_i_2__3 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[20]),
        .I2(STALL_EN),
        .I3(IF_PC2[20]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[20] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[20]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000E2)) 
    \Q[20]_i_3 
       (.I0(\Q[20]_i_11__1_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[23]_i_15_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [7]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [6]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [19]));
  LUT6 #(
    .INIT(64'hFCFFFCDDFCCCFCDD)) 
    \Q[20]_i_3__0 
       (.I0(\Q[20]_i_5__0_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [18]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[20]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFFFBFAF)) 
    \Q[20]_i_3__1 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(\custom_alu/fp2int/INT0 [15]),
        .I2(EX_CUSTOM_ALU_SEL[27]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/fp2int/p_0_in [15]),
        .O(\Q[20]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[20]_i_3__2 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(data1[5]),
        .O(\Q[20]_i_3__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[20]_i_3__3 
       (.I0(EX_MEM_Q[39]),
        .I1(EX_MEM_Q[37]),
        .O(MEM_D_MEM_ALU_FINAL1));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[20]_i_3__4 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[19]),
        .I2(STALL_EN),
        .I3(IF_PC2[19]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[19] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[20]_i_3__4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000E2)) 
    \Q[20]_i_4 
       (.I0(\Q[20]_i_12__1_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[20]_i_11__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [7]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [6]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [18]));
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT4 #(
    .INIT(16'hBBFB)) 
    \Q[20]_i_4__0 
       (.I0(\custom_alu/fp32_add/sel0 [23]),
        .I1(\custom_alu/fp32_add/sel0 [24]),
        .I2(\custom_alu/fp32_add/sel0 [22]),
        .I3(\custom_alu/fp32_add/sel0 [19]),
        .O(\Q[20]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h4FFF4F4F44444444)) 
    \Q[20]_i_4__1 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [15]),
        .I2(\Q[20]_i_7__0_n_0 ),
        .I3(\Q[20]_i_8__0_n_0 ),
        .I4(\Q[26]_i_7_n_0 ),
        .I5(\Q[30]_i_5_n_0 ),
        .O(\Q[20]_i_4__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \Q[20]_i_4__2 
       (.I0(MEM_LOAD_SEL[5]),
        .I1(MEM_LOAD_SEL[6]),
        .O(\Q[20]_i_4__2_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[20]_i_4__3 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[18]),
        .I2(STALL_EN),
        .I3(IF_PC2[18]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[18] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[20]_i_4__3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000E2)) 
    \Q[20]_i_5 
       (.I0(\Q[20]_i_13__1_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[20]_i_12__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [7]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [6]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [17]));
  LUT6 #(
    .INIT(64'h00000000FFFFEEFE)) 
    \Q[20]_i_5__0 
       (.I0(\custom_alu/fp32_add/sel0 [19]),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [17]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\Q[20]_i_6__0_n_0 ),
        .I5(\Q[20]_i_7_n_0 ),
        .O(\Q[20]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    \Q[20]_i_5__1 
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__2_i_7_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__2_i_5_n_0),
        .O(\custom_alu/fp2int/p_0_in [15]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[20]_i_5__2 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[17]),
        .I2(STALL_EN),
        .I3(IF_PC2[17]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[17] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[20]_i_5__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000E2)) 
    \Q[20]_i_6 
       (.I0(\Q[20]_i_14__1_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[20]_i_13__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [7]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [6]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [16]));
  LUT6 #(
    .INIT(64'h0030023203330232)) 
    \Q[20]_i_6__0 
       (.I0(\Q[20]_i_8_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [16]),
        .I3(\custom_alu/fp32_add/sel0 [13]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[20]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT4 #(
    .INIT(16'hB888)) 
    \Q[20]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [16]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [15]),
        .I3(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000553FFFFF553F)) 
    \Q[20]_i_7__0 
       (.I0(\Q[31]_i_14__0_n_0 ),
        .I1(\Q[31]_i_11__0_n_0 ),
        .I2(\Q[35]_i_16_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .I5(\Q[31]_i_13__0_n_0 ),
        .O(\Q[20]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h002AAA2A)) 
    \Q[20]_i_8 
       (.I0(\Q[20]_i_9_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [13]),
        .I2(\custom_alu/fp32_add/sel0 [10]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAAA2)) 
    \Q[20]_i_8__0 
       (.I0(\Q[30]_i_8_n_0 ),
        .I1(\Q[30]_i_9__0_n_0 ),
        .I2(\Q[27]_i_13_n_0 ),
        .I3(\Q[20]_i_13__0_n_0 ),
        .I4(\Q[20]_i_14_n_0 ),
        .I5(\Q[30]_i_11__0_n_0 ),
        .O(\Q[20]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \Q[20]_i_9 
       (.I0(\Q[20]_i_10_n_0 ),
        .I1(\Q[20]_i_11_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [12]),
        .I3(\custom_alu/fp32_add/sel0 [9]),
        .I4(\custom_alu/fp32_add/sel0 [13]),
        .I5(\custom_alu/fp32_add/sel0 [14]),
        .O(\Q[20]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[20]_i_9__0 
       (.I0(exponent_carry_i_10_n_7),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_11_n_4),
        .O(\Q[20]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[21]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [21]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [20]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [21]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF02F2)) 
    \Q[21]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [4]),
        .I2(\custom_alu/fp32_add/sel0 [7]),
        .I3(\custom_alu/fp32_add/sel0 [5]),
        .I4(\custom_alu/fp32_add/sel0 [8]),
        .I5(\custom_alu/fp32_add/sel0 [9]),
        .O(\Q[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEFEAFFFAEFEFFFFF)) 
    \Q[21]_i_10__0 
       (.I0(\Q[31]_i_14__0_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [20]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN1[20]),
        .I4(\custom_alu/int2fp/INT_VAL0 [19]),
        .I5(ALU_DIN1[19]),
        .O(\Q[21]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000007577)) 
    \Q[21]_i_11 
       (.I0(\custom_alu/fp32_add/sel0 [3]),
        .I1(\custom_alu/fp32_add/sel0 [5]),
        .I2(\custom_alu/fp32_add/sel0 [4]),
        .I3(\custom_alu/fp32_add/sel0 [1]),
        .I4(\Q[21]_i_12_n_0 ),
        .I5(\Q[21]_i_13_n_0 ),
        .O(\Q[21]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8888888B888)) 
    \Q[21]_i_11__0 
       (.I0(\Q[17]_i_11__0_n_0 ),
        .I1(\Q[31]_i_14__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(ALU_DIN1[13]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [13]),
        .O(\Q[21]_i_11__0_n_0 ));
  LUT5 #(
    .INIT(32'h44440040)) 
    \Q[21]_i_12 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [2]),
        .I2(\custom_alu/fp32_add/sel0 [0]),
        .I3(\custom_alu/fp32_add/sel0 [3]),
        .I4(\custom_alu/fp32_add/sel0 [4]),
        .O(\Q[21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8B8B88B888888)) 
    \Q[21]_i_12__0 
       (.I0(\Q[69]_i_16_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[17]_i_14_n_0 ),
        .I4(\Q[31]_i_13__0_n_0 ),
        .I5(\Q[17]_i_10__0_n_0 ),
        .O(\Q[21]_i_12__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \Q[21]_i_13 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [7]),
        .O(\Q[21]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAEFF00)) 
    \Q[21]_i_1__0 
       (.I0(\Q[21]_i_2_n_0 ),
        .I1(\Q[21]_i_3_n_0 ),
        .I2(\Q[21]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[22] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [21]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[21]_i_1__1 
       (.I0(\Q[21]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[6]),
        .I3(data1[6]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[6]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[21]_i_1__2 
       (.I0(\Q[21]_i_2__0_n_0 ),
        .I1(\Q[21]_i_3__0_n_0 ),
        .I2(\Q[21]_i_4__0_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[16]),
        .O(data0[16]));
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT5 #(
    .INIT(32'hFFFFEAEE)) 
    \Q[21]_i_1__3 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[21]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(\Q[21]_i_2__2_n_0 ),
        .O(data1[16]));
  LUT4 #(
    .INIT(16'h8F80)) 
    \Q[21]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [21]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [24]),
        .I3(\custom_alu/fp32_add/data23 [21]),
        .O(\Q[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[21]_i_2__0 
       (.I0(\custom_alu/MULT [16]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [48]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [16]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[21]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[21]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[6]),
        .I2(CRF_RD2_IBUF[6]),
        .I3(RF_RD2_IBUF[6]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[21]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT5 #(
    .INIT(32'h0000A280)) 
    \Q[21]_i_2__2 
       (.I0(\Q[21]_i_3__1_n_0 ),
        .I1(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I2(D_MEM_DOUT_IBUF[24]),
        .I3(D_MEM_DOUT_IBUF[16]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .O(\Q[21]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFFCDDFCCCFCDD)) 
    \Q[21]_i_3 
       (.I0(\Q[21]_i_5_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [19]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [20]),
        .I5(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[21]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hBFFFBFAF)) 
    \Q[21]_i_3__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(\custom_alu/fp2int/INT0 [16]),
        .I2(EX_CUSTOM_ALU_SEL[27]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/fp2int/p_0_in [16]),
        .O(\Q[21]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \Q[21]_i_3__1 
       (.I0(MEM_LOAD_SEL[5]),
        .I1(MEM_LOAD_SEL[6]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(MEM_LOAD_SEL[2]),
        .I5(MEM_LOAD_SEL[1]),
        .O(\Q[21]_i_3__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT4 #(
    .INIT(16'hBBFB)) 
    \Q[21]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [23]),
        .I1(\custom_alu/fp32_add/sel0 [24]),
        .I2(\custom_alu/fp32_add/sel0 [22]),
        .I3(\custom_alu/fp32_add/sel0 [20]),
        .O(\Q[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF44F444444444)) 
    \Q[21]_i_4__0 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [16]),
        .I2(\Q[26]_i_7_n_0 ),
        .I3(\Q[21]_i_6__0_n_0 ),
        .I4(\Q[21]_i_7__0_n_0 ),
        .I5(\Q[30]_i_5_n_0 ),
        .O(\Q[21]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h10DC13DC13DF13DF)) 
    \Q[21]_i_5 
       (.I0(\custom_alu/fp32_add/sel0 [16]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [18]),
        .I3(\custom_alu/fp32_add/sel0 [17]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\Q[21]_i_6_n_0 ),
        .O(\Q[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    \Q[21]_i_5__0 
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__2_i_5_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__2_i_6_n_0),
        .O(\custom_alu/fp2int/p_0_in [16]));
  LUT6 #(
    .INIT(64'hFFCFFDCDFCCCFDCD)) 
    \Q[21]_i_6 
       (.I0(\Q[21]_i_7_n_0 ),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [16]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\custom_alu/fp32_add/sel0 [13]),
        .O(\Q[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0DDD00000DDD0DDD)) 
    \Q[21]_i_6__0 
       (.I0(\Q[21]_i_8__0_n_0 ),
        .I1(\Q[21]_i_9__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[35]_i_17_n_0 ),
        .I4(\Q[31]_i_7_n_0 ),
        .I5(\Q[31]_i_6_n_0 ),
        .O(\Q[21]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'h553F5530)) 
    \Q[21]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [12]),
        .I1(\custom_alu/fp32_add/sel0 [11]),
        .I2(\custom_alu/fp32_add/sel0 [13]),
        .I3(\custom_alu/fp32_add/sel0 [14]),
        .I4(\Q[21]_i_8_n_0 ),
        .O(\Q[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[21]_i_7__0 
       (.I0(\Q[28]_i_20_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[31]_i_13__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[21]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFF1D1D3F0C)) 
    \Q[21]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [11]),
        .I2(\custom_alu/fp32_add/sel0 [9]),
        .I3(\Q[21]_i_9_n_0 ),
        .I4(\custom_alu/fp32_add/sel0 [10]),
        .I5(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[21]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00F2)) 
    \Q[21]_i_8__0 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\Q[21]_i_10__0_n_0 ),
        .I2(\Q[21]_i_11__0_n_0 ),
        .I3(\Q[67]_i_12_n_0 ),
        .I4(\Q[21]_i_12__0_n_0 ),
        .I5(\Q[29]_i_7_n_0 ),
        .O(\Q[21]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000EEEEEEE0EEE)) 
    \Q[21]_i_9 
       (.I0(\Q[21]_i_10_n_0 ),
        .I1(\Q[21]_i_11_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [8]),
        .I3(\custom_alu/fp32_add/sel0 [6]),
        .I4(\custom_alu/fp32_add/sel0 [9]),
        .I5(\custom_alu/fp32_add/sel0 [7]),
        .O(\Q[21]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \Q[21]_i_9__0 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[31]_i_10__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[21]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[22]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [22]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [21]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [22]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[22]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[22]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF000E000F0000000)) 
    \Q[22]_i_10__0 
       (.I0(\Q[22]_i_16__0_n_0 ),
        .I1(\Q[67]_i_12_n_0 ),
        .I2(\Q[27]_i_13_n_0 ),
        .I3(\Q[22]_i_17_n_0 ),
        .I4(\Q[9]_i_11_n_0 ),
        .I5(\Q[22]_i_18__0_n_0 ),
        .O(\Q[22]_i_10__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[22]_i_11 
       (.I0(\custom_alu/fp32_add/sel0 [17]),
        .O(\Q[22]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    \Q[22]_i_11__0 
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__2_i_6_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__3_i_8_n_0),
        .O(\custom_alu/fp2int/p_0_in [17]));
  LUT6 #(
    .INIT(64'h0000FFFF0F0F3437)) 
    \Q[22]_i_12 
       (.I0(\custom_alu/fp32_add/sel0 [14]),
        .I1(\custom_alu/fp32_add/sel0 [15]),
        .I2(\custom_alu/fp32_add/sel0 [16]),
        .I3(\Q[22]_i_13_n_0 ),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .I5(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[22]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFF47444744)) 
    \Q[22]_i_12__0 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[17]_i_11__0_n_0 ),
        .I2(\Q[35]_i_26_n_0 ),
        .I3(\Q[28]_i_18_n_0 ),
        .I4(\Q[35]_i_22_n_0 ),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[22]_i_12__0_n_0 ));
  LUT5 #(
    .INIT(32'hFA03FA00)) 
    \Q[22]_i_13 
       (.I0(\custom_alu/fp32_add/sel0 [12]),
        .I1(\Q[22]_i_14_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [14]),
        .I3(\custom_alu/fp32_add/sel0 [13]),
        .I4(\Q[22]_i_15_n_0 ),
        .O(\Q[22]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[22]_i_13__0 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_20_n_0 ),
        .I2(\Q[35]_i_28_n_0 ),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[22]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00F1)) 
    \Q[22]_i_14 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\Q[22]_i_16_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [10]),
        .I3(\custom_alu/fp32_add/sel0 [9]),
        .I4(\custom_alu/fp32_add/sel0 [12]),
        .I5(\custom_alu/fp32_add/sel0 [11]),
        .O(\Q[22]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h0000F808)) 
    \Q[22]_i_14__0 
       (.I0(\Q[47]_i_9_n_0 ),
        .I1(\Q[35]_i_26_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[35]_i_32_n_0 ),
        .I4(\Q[35]_i_22_n_0 ),
        .O(\Q[22]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FF0E)) 
    \Q[22]_i_15 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\Q[22]_i_17__0_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [9]),
        .I3(\custom_alu/fp32_add/sel0 [8]),
        .I4(\custom_alu/fp32_add/sel0 [11]),
        .I5(\Q[22]_i_18_n_0 ),
        .O(\Q[22]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF000800000008)) 
    \Q[22]_i_15__0 
       (.I0(ALU_DIN1[0]),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[35]_i_22_n_0 ),
        .I5(\Q[29]_i_18__0_n_0 ),
        .O(\Q[22]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00F2)) 
    \Q[22]_i_16 
       (.I0(\custom_alu/fp32_add/sel0 [1]),
        .I1(\custom_alu/fp32_add/sel0 [4]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [6]),
        .I4(\custom_alu/fp32_add/sel0 [5]),
        .I5(\custom_alu/fp32_add/sel0 [8]),
        .O(\Q[22]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000F77FFFF0F77)) 
    \Q[22]_i_16__0 
       (.I0(\Q[28]_i_18_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[31]_i_11__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[22]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000535FFFFF535F)) 
    \Q[22]_i_17 
       (.I0(\Q[31]_i_11__0_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[23]_i_13__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[31]_i_14__0_n_0 ),
        .O(\Q[22]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h4544454545444544)) 
    \Q[22]_i_17__0 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [4]),
        .I2(\custom_alu/fp32_add/sel0 [5]),
        .I3(\custom_alu/fp32_add/sel0 [2]),
        .I4(\custom_alu/fp32_add/sel0 [3]),
        .I5(\custom_alu/fp32_add/sel0 [0]),
        .O(\Q[22]_i_17__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \Q[22]_i_18 
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .O(\Q[22]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h5530553F553F553F)) 
    \Q[22]_i_18__0 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[29]_i_10_n_0 ),
        .I4(\Q[17]_i_10__0_n_0 ),
        .I5(\Q[31]_i_13__0_n_0 ),
        .O(\Q[22]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F2F2FF00)) 
    \Q[22]_i_1__0 
       (.I0(\custom_alu/fp32_add/data23 [22]),
        .I1(\custom_alu/fp32_add/sel0 [24]),
        .I2(\Q[22]_i_3_n_0 ),
        .I3(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[23] ),
        .I4(\Q[30]_i_2__1_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [22]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[22]_i_1__1 
       (.I0(\Q[22]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[7]),
        .I3(data1[7]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[7]));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[22]_i_1__2 
       (.I0(\Q[22]_i_2_n_0 ),
        .I1(\Q[22]_i_3__0_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[17]),
        .O(data0[17]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[22]_i_1__3 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[22]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[17]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[17]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[22]_i_2 
       (.I0(\custom_alu/MULT [17]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [49]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(\custom_alu/Q [17]),
        .O(\Q[22]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[22]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[7]),
        .I2(CRF_RD2_IBUF[7]),
        .I3(RF_RD2_IBUF[7]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[22]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FC000000F800)) 
    \Q[22]_i_3 
       (.I0(\custom_alu/fp32_add/sel0 [20]),
        .I1(\custom_alu/fp32_add/sel0 [21]),
        .I2(\Q[22]_i_7_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\custom_alu/fp32_add/sel0 [23]),
        .I5(\custom_alu/fp32_add/sel0 [22]),
        .O(\Q[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h7500000075007500)) 
    \Q[22]_i_3__0 
       (.I0(\Q[30]_i_5_n_0 ),
        .I1(\Q[22]_i_4_n_0 ),
        .I2(\Q[22]_i_5__0_n_0 ),
        .I3(\Q[22]_i_6__0_n_0 ),
        .I4(\Q[65]_i_5_n_0 ),
        .I5(\custom_alu/fp32_mult/product_mantissa [17]),
        .O(\Q[22]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF0D0000)) 
    \Q[22]_i_4 
       (.I0(\Q[22]_i_7__0_n_0 ),
        .I1(\Q[22]_i_8__0_n_0 ),
        .I2(\Q[22]_i_9__0_n_0 ),
        .I3(\Q[27]_i_13_n_0 ),
        .I4(\Q[26]_i_7_n_0 ),
        .I5(\Q[22]_i_10__0_n_0 ),
        .O(\Q[22]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[22]_i_5 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .O(\Q[22]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000553FFFFF553F)) 
    \Q[22]_i_5__0 
       (.I0(\Q[28]_i_20_n_0 ),
        .I1(\Q[31]_i_13__0_n_0 ),
        .I2(\Q[35]_i_16_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .I5(\Q[29]_i_10_n_0 ),
        .O(\Q[22]_i_5__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[22]_i_6 
       (.I0(\custom_alu/fp32_add/sel0 [21]),
        .O(\Q[22]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBFFFBFAF)) 
    \Q[22]_i_6__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(\custom_alu/fp2int/INT0 [17]),
        .I2(EX_CUSTOM_ALU_SEL[27]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/fp2int/p_0_in [17]),
        .O(\Q[22]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h1100110110001001)) 
    \Q[22]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .I1(\custom_alu/fp32_add/sel0 [21]),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [19]),
        .I4(\Q[22]_i_12_n_0 ),
        .I5(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000003000355)) 
    \Q[22]_i_7__0 
       (.I0(ALU_DIN1[17]),
        .I1(\custom_alu/int2fp/INT_VAL0 [17]),
        .I2(\custom_alu/int2fp/INT_VAL0 [16]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN1[16]),
        .I5(\Q[28]_i_11_n_0 ),
        .O(\Q[22]_i_7__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[22]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [20]),
        .O(\Q[22]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5555555055554444)) 
    \Q[22]_i_8__0 
       (.I0(\Q[22]_i_12__0_n_0 ),
        .I1(\Q[22]_i_13__0_n_0 ),
        .I2(\Q[22]_i_14__0_n_0 ),
        .I3(\Q[22]_i_15__0_n_0 ),
        .I4(\Q[26]_i_20_n_0 ),
        .I5(\Q[26]_i_23_n_0 ),
        .O(\Q[22]_i_8__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[22]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [19]),
        .O(\Q[22]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0002FF0200F2FFF2)) 
    \Q[22]_i_9__0 
       (.I0(\Q[17]_i_10__0_n_0 ),
        .I1(\Q[35]_i_21_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[35]_i_20_n_0 ),
        .I5(\Q[35]_i_19_n_0 ),
        .O(\Q[22]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h0B08)) 
    \Q[23]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [23]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\Q[30]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/significand_add0 [22]),
        .O(\custom_alu/fp32_add/p_1_out [23]));
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \Q[23]_i_11 
       (.I0(\Q[23]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .O(\Q[23]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000005404)) 
    \Q[23]_i_12 
       (.I0(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I1(ALU_DIN2[22]),
        .I2(\custom_alu/fp32_add/op_a2 ),
        .I3(ALU_DIN1[22]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [2]),
        .O(\Q[23]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \Q[23]_i_13 
       (.I0(\custom_alu/fp32_add/p_1_in__0 [6]),
        .I1(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [7]),
        .O(\Q[23]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[23]_i_13__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [25]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[151]),
        .I5(EX_RF_RD1[25]),
        .O(\Q[23]_i_13__0_n_0 ));
  LUT5 #(
    .INIT(32'h88888B88)) 
    \Q[23]_i_14 
       (.I0(\Q[23]_i_11_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I3(\Q[23]_i_19_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [2]),
        .O(\Q[23]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h10131010DCDFDCDC)) 
    \Q[23]_i_14__0 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\Q[28]_i_11_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[17]_i_10__0_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[23]_i_14__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000B08)) 
    \Q[23]_i_15 
       (.I0(\Q[23]_i_20_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I3(\Q[23]_i_21_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [2]),
        .O(\Q[23]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFD5DFD5DFD5DF)) 
    \Q[23]_i_15__0 
       (.I0(\Q[69]_i_20_n_0 ),
        .I1(\Q[17]_i_15_n_0 ),
        .I2(\Q[35]_i_22_n_0 ),
        .I3(\Q[23]_i_16__0_n_0 ),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[35]_i_27_n_0 ),
        .O(\Q[23]_i_15__0_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[23]_i_16 
       (.I0(ID_EX_Q[100]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[21]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[21]),
        .O(\Q[23]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0074FF74)) 
    \Q[23]_i_16__0 
       (.I0(\Q[47]_i_9_n_0 ),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[23]_i_17__0_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[35]_i_32_n_0 ),
        .I5(\Q[35]_i_27_n_0 ),
        .O(\Q[23]_i_16__0_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[23]_i_17 
       (.I0(ID_EX_Q[99]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[20]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[20]),
        .O(\Q[23]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \Q[23]_i_17__0 
       (.I0(ALU_DIN1[0]),
        .I1(EX_RF_RD1[5]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[131]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\custom_alu/int2fp/INT_VAL0 [5]),
        .O(\Q[23]_i_17__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \Q[23]_i_18 
       (.I0(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I1(\Q[23]_i_22_n_0 ),
        .O(\Q[23]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[23]_i_19 
       (.I0(EX_RF_RD2[21]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[100]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[21]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[23]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[23]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[24] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [0]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [23]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[23]_i_1__1 
       (.I0(\Q[23]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[8]),
        .I3(data1[8]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[8]));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[23]_i_1__2 
       (.I0(\Q[23]_i_2_n_0 ),
        .I1(\Q[23]_i_3__0_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[18]),
        .O(data0[18]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[23]_i_1__3 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[23]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[18]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[23]_i_1__4 
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[23]),
        .O(ALU_DIN2[23]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[23]_i_2 
       (.I0(\custom_alu/MULT [18]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [50]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(\custom_alu/Q [18]),
        .O(\Q[23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[23]_i_20 
       (.I0(EX_RF_RD2[22]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[101]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[22]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[23]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[23]_i_21 
       (.I0(EX_RF_RD2[20]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[99]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[20]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[23]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \Q[23]_i_22 
       (.I0(\custom_alu/fp32_add/p_0_in2_in [5]),
        .I1(\custom_alu/fp32_add/p_0_in2_in [6]),
        .I2(\custom_alu/fp32_add/p_0_in2_in [1]),
        .I3(\custom_alu/fp32_add/p_0_in2_in [2]),
        .I4(\Q[23]_i_23_n_0 ),
        .O(\Q[23]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFEFEFE)) 
    \Q[23]_i_23 
       (.I0(\custom_alu/fp32_add/p_0_in2_in [3]),
        .I1(\custom_alu/fp32_add/p_0_in2_in [0]),
        .I2(\custom_alu/fp32_add/p_0_in2_in [4]),
        .I3(ALU_DIN1[30]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[30]),
        .O(\Q[23]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[23]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[8]),
        .I2(CRF_RD2_IBUF[8]),
        .I3(RF_RD2_IBUF[8]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[23]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \Q[23]_i_3 
       (.I0(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I1(\Q[23]_i_11_n_0 ),
        .I2(\custom_alu/fp32_add/p_1_in__0 [6]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [7]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [0]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [23]));
  LUT6 #(
    .INIT(64'h000000000BBB0B0B)) 
    \Q[23]_i_3__0 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [18]),
        .I2(\Q[30]_i_5_n_0 ),
        .I3(\Q[23]_i_6__0_n_0 ),
        .I4(\Q[23]_i_7_n_0 ),
        .I5(\Q[65]_i_8_n_0 ),
        .O(\Q[23]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h00005404)) 
    \Q[23]_i_4 
       (.I0(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I1(\Q[23]_i_12_n_0 ),
        .I2(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I3(\Q[23]_i_11_n_0 ),
        .I4(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [22]));
  LUT5 #(
    .INIT(32'h00002E22)) 
    \Q[23]_i_5 
       (.I0(\Q[23]_i_14_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I3(\Q[23]_i_12_n_0 ),
        .I4(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [21]));
  LUT6 #(
    .INIT(64'h00000000000000E2)) 
    \Q[23]_i_6 
       (.I0(\Q[23]_i_15_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[23]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [7]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [6]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [20]));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[23]_i_6__0 
       (.I0(\Q[23]_i_13__0_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[29]_i_10_n_0 ),
        .I4(\Q[28]_i_20_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFB0000FFFFFFFF)) 
    \Q[23]_i_7 
       (.I0(\Q[23]_i_14__0_n_0 ),
        .I1(\Q[23]_i_15__0_n_0 ),
        .I2(\Q[27]_i_13_n_0 ),
        .I3(\Q[65]_i_14_n_0 ),
        .I4(\Q[65]_i_15_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFE)) 
    \Q[23]_i_7__0 
       (.I0(\Q[87]_i_12_n_0 ),
        .I1(\custom_alu/fp32_add/p_0_in [2]),
        .I2(\custom_alu/fp32_add/p_0_in [3]),
        .I3(\custom_alu/fp32_add/p_0_in [1]),
        .I4(\custom_alu/fp32_add/p_0_in [0]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [23]),
        .O(\Q[23]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'hE21DE2E2)) 
    \Q[24]_i_1 
       (.I0(ALU_DIN1[23]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN2[23]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .I4(\custom_alu/fp32_add/significand_add0 [24]),
        .O(\custom_alu/fp32_add/p_1_out [24]));
  LUT6 #(
    .INIT(64'hAAABAAABAAABAAAA)) 
    \Q[24]_i_10 
       (.I0(\Q[24]_i_15_n_0 ),
        .I1(\Q[69]_i_20_n_0 ),
        .I2(\Q[27]_i_13_n_0 ),
        .I3(\Q[24]_i_16_n_0 ),
        .I4(\Q[24]_i_17_n_0 ),
        .I5(\Q[24]_i_18_n_0 ),
        .O(\Q[24]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[24]_i_11 
       (.I0(\Q[17]_i_10__0_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[17]_i_14_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[17]_i_11__0_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[24]_i_12 
       (.I0(\Q[35]_i_28_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[35]_i_29_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[35]_i_26_n_0 ),
        .O(\Q[24]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h4447474774777777)) 
    \Q[24]_i_13 
       (.I0(\Q[35]_i_21_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[31]_i_13__0_n_0 ),
        .I4(\Q[35]_i_27_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[24]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \Q[24]_i_14 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[35]_i_20_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \Q[24]_i_15 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(EX_RF_RD1[13]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[139]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [13]),
        .O(\Q[24]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \Q[24]_i_16 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(EX_RF_RD1[4]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[130]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [4]),
        .O(\Q[24]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h3033302230003022)) 
    \Q[24]_i_17 
       (.I0(\Q[24]_i_19_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[35]_i_32_n_0 ),
        .I3(\Q[17]_i_10__0_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[47]_i_9_n_0 ),
        .O(\Q[24]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hEFEAAFAAEAEAAAAA)) 
    \Q[24]_i_18 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [17]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN1[17]),
        .I4(\custom_alu/int2fp/INT_VAL0 [3]),
        .I5(ALU_DIN1[3]),
        .O(\Q[24]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \Q[24]_i_19 
       (.I0(EX_RF_RD1[14]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[140]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [14]),
        .I5(ALU_DIN1[0]),
        .O(\Q[24]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[24]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[25] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [1]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [24]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[24]_i_1__1 
       (.I0(\Q[24]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[9]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[9]),
        .I5(\Q[24]_i_4__0_n_0 ),
        .O(ID_RD2_FORWARDED[9]));
  LUT6 #(
    .INIT(64'hBBBAFFFFBBBA0000)) 
    \Q[24]_i_1__2 
       (.I0(\Q[24]_i_2_n_0 ),
        .I1(\Q[24]_i_3__1_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\Q[24]_i_4_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[19]),
        .O(data0[19]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[24]_i_1__3 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[24]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[19]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[19]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[24]_i_1__4 
       (.I0(ID_EX_Q[103]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[24]),
        .O(ALU_DIN2[24]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[24]_i_2 
       (.I0(\custom_alu/MULT [19]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [51]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [19]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[24]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[9]),
        .I2(CRF_RD2_IBUF[9]),
        .I3(RF_RD2_IBUF[9]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[24]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[24]_i_2__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[24]),
        .I2(STALL_EN),
        .I3(IF_PC2[24]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[24] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[24]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hBBBFBBBBAAAAAAAA)) 
    \Q[24]_i_3 
       (.I0(\Q[14]_i_2__0_n_0 ),
        .I1(\Q[24]_i_5__1_n_0 ),
        .I2(\Q[24]_i_6__0_n_0 ),
        .I3(\Q[24]_i_7__0_n_0 ),
        .I4(\Q[24]_i_8__0_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[9]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[24]_i_3__0 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[23]),
        .I2(STALL_EN),
        .I3(IF_PC2[23]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[23] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[24]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    \Q[24]_i_3__1 
       (.I0(\custom_alu/fp32_mult/product_mantissa [19]),
        .I1(\Q[25]_i_5_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(EX_CUSTOM_ALU_SEL[31]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(EX_CUSTOM_ALU_SEL[30]),
        .O(\Q[24]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hF0220022F022FF22)) 
    \Q[24]_i_4 
       (.I0(EX_CUSTOM_ALU_SEL[26]),
        .I1(\Q[24]_i_5_n_0 ),
        .I2(\custom_alu/fp2int/INT0 [19]),
        .I3(EX_CUSTOM_ALU_SEL[27]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\custom_alu/fp2int/p_0_in [19]),
        .O(\Q[24]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \Q[24]_i_4__0 
       (.I0(DIN2_FORWARD[0]),
        .I1(DIN2_FORWARD[1]),
        .I2(data1[9]),
        .O(\Q[24]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[24]_i_4__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[22]),
        .I2(STALL_EN),
        .I3(IF_PC2[22]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[22] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[24]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555DDFD)) 
    \Q[24]_i_5 
       (.I0(\Q[26]_i_7_n_0 ),
        .I1(\Q[24]_i_7_n_0 ),
        .I2(\Q[35]_i_17_n_0 ),
        .I3(\Q[28]_i_20_n_0 ),
        .I4(\Q[24]_i_8_n_0 ),
        .I5(\Q[66]_i_7_n_0 ),
        .O(\Q[24]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[24]_i_5__0 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[21]),
        .I2(STALL_EN),
        .I3(IF_PC2[21]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[21] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[24]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFEFFFFF)) 
    \Q[24]_i_5__1 
       (.I0(\Q[69]_i_13_n_0 ),
        .I1(\Q[69]_i_14_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .I4(\custom_alu/fp32_mult/product_mantissa [9]),
        .O(\Q[24]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    \Q[24]_i_6 
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__3_i_7_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__3_i_5_n_0),
        .O(\custom_alu/fp2int/p_0_in [19]));
  LUT6 #(
    .INIT(64'h0000115155555555)) 
    \Q[24]_i_6__0 
       (.I0(EX_CUSTOM_ALU_SEL[27]),
        .I1(\Q[26]_i_7_n_0 ),
        .I2(\Q[24]_i_9_n_0 ),
        .I3(\Q[24]_i_10_n_0 ),
        .I4(\Q[24]_i_11_n_0 ),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[24]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000022202220222)) 
    \Q[24]_i_7 
       (.I0(\Q[66]_i_18_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[31]_i_13__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[28]_i_21_n_0 ),
        .O(\Q[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[24]_i_7__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [9]),
        .O(\Q[24]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h000055FD)) 
    \Q[24]_i_8 
       (.I0(\Q[22]_i_7__0_n_0 ),
        .I1(\Q[66]_i_13_n_0 ),
        .I2(\Q[24]_i_9__0_n_0 ),
        .I3(\Q[66]_i_11_n_0 ),
        .I4(\Q[66]_i_9_n_0 ),
        .O(\Q[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0047FFFFFFFF)) 
    \Q[24]_i_8__0 
       (.I0(INT0_carry__1_i_14_n_0),
        .I1(ALU_DIN1[23]),
        .I2(INT0_carry__0_i_6_n_0),
        .I3(INT0_carry_i_6_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[24]_i_8__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5400)) 
    \Q[24]_i_9 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[24]_i_12_n_0 ),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[24]_i_13_n_0 ),
        .I4(\Q[24]_i_14_n_0 ),
        .O(\Q[24]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[24]_i_9__0 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[35]_i_20_n_0 ),
        .I2(\Q[35]_i_26_n_0 ),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[35]_i_29_n_0 ),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[24]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'hA6AAA6A6A6AAAAAA)) 
    \Q[25]_i_1 
       (.I0(\custom_alu/fp32_add/p_0_in [1]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\Q[30]_i_4__0_n_0 ),
        .I3(ALU_DIN2[23]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN1[23]),
        .O(\custom_alu/fp32_add/p_1_out [25]));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[25]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[26] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [2]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [25]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[25]_i_1__1 
       (.I0(\Q[25]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[10]),
        .I3(data1[10]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[10]));
  LUT6 #(
    .INIT(64'hBBBAFFFFBBBA0000)) 
    \Q[25]_i_1__2 
       (.I0(\Q[25]_i_2_n_0 ),
        .I1(\Q[25]_i_3_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\Q[25]_i_4_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[20]),
        .O(data0[20]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[25]_i_1__3 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[25]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[20]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[25]_i_1__4 
       (.I0(ID_EX_Q[104]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[25]),
        .O(ALU_DIN2[25]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[25]_i_2 
       (.I0(\custom_alu/MULT [20]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [52]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [20]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[25]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[10]),
        .I2(CRF_RD2_IBUF[10]),
        .I3(RF_RD2_IBUF[10]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[25]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    \Q[25]_i_3 
       (.I0(\custom_alu/fp32_mult/product_mantissa [20]),
        .I1(\Q[25]_i_5_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(EX_CUSTOM_ALU_SEL[31]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(EX_CUSTOM_ALU_SEL[30]),
        .O(\Q[25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0220022F022FF22)) 
    \Q[25]_i_4 
       (.I0(EX_CUSTOM_ALU_SEL[26]),
        .I1(\Q[25]_i_6_n_0 ),
        .I2(\custom_alu/fp2int/INT0 [20]),
        .I3(EX_CUSTOM_ALU_SEL[27]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/fp2int/p_0_in [20]),
        .O(\Q[25]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \Q[25]_i_5 
       (.I0(\Q[69]_i_14_n_0 ),
        .I1(\Q[69]_i_13_n_0 ),
        .I2(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .O(\Q[25]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h77773333777700F0)) 
    \Q[25]_i_6 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(\Q[25]_i_8_n_0 ),
        .I2(\Q[67]_i_8_n_0 ),
        .I3(\Q[67]_i_9__0_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .I5(\Q[26]_i_15__0_n_0 ),
        .O(\Q[25]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEAEAEFEFEAEFE)) 
    \Q[25]_i_7 
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__3_i_5_n_0),
        .I2(ALU_DIN1[23]),
        .I3(ALU_DIN1[24]),
        .I4(INT0_carry__3_i_6_n_0),
        .I5(ALU_DIN1[21]),
        .O(\custom_alu/fp2int/p_0_in [20]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \Q[25]_i_8 
       (.I0(\Q[28]_i_7_n_0 ),
        .I1(\Q[23]_i_13__0_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[28]_i_12_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .O(\Q[25]_i_8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[26]_i_1 
       (.I0(\Q[27]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[28]),
        .O(CUSTOM_ALU_SEL[26]));
  LUT6 #(
    .INIT(64'hBABFBABABABFBEBE)) 
    \Q[26]_i_10 
       (.I0(\Q[27]_i_13_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[28]_i_11_n_0 ),
        .I3(\Q[17]_i_14_n_0 ),
        .I4(\Q[69]_i_16_n_0 ),
        .I5(\Q[17]_i_11__0_n_0 ),
        .O(\Q[26]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000AB)) 
    \Q[26]_i_10__0 
       (.I0(\Q[26]_i_16__0_n_0 ),
        .I1(\Q[35]_i_23_n_0 ),
        .I2(\Q[26]_i_17_n_0 ),
        .I3(\Q[26]_i_18_n_0 ),
        .I4(\Q[27]_i_13_n_0 ),
        .I5(\Q[69]_i_20_n_0 ),
        .O(\Q[26]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'hBABABABEBFBABFBE)) 
    \Q[26]_i_11 
       (.I0(\Q[26]_i_20_n_0 ),
        .I1(\Q[35]_i_21_n_0 ),
        .I2(\Q[35]_i_20_n_0 ),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[35]_i_27_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[26]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[26]_i_11__0 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[69]_i_16_n_0 ),
        .I4(\Q[17]_i_10__0_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[26]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \Q[26]_i_12 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(EX_RF_RD1[15]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[141]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\custom_alu/int2fp/INT_VAL0 [15]),
        .O(\Q[26]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h88A8888800000000)) 
    \Q[26]_i_12__0 
       (.I0(\Q[26]_i_21_n_0 ),
        .I1(\Q[26]_i_22_n_0 ),
        .I2(ALU_DIN1[0]),
        .I3(\Q[29]_i_18__0_n_0 ),
        .I4(\Q[35]_i_32_n_0 ),
        .I5(\Q[69]_i_22_n_0 ),
        .O(\Q[26]_i_12__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \Q[26]_i_13 
       (.I0(\Q[28]_i_21_n_0 ),
        .I1(\Q[28]_i_18_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[17]_i_11__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[26]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCF808FFFFFFFF)) 
    \Q[26]_i_13__0 
       (.I0(\Q[35]_i_28_n_0 ),
        .I1(\Q[35]_i_26_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[35]_i_29_n_0 ),
        .I4(\Q[35]_i_22_n_0 ),
        .I5(\Q[26]_i_23_n_0 ),
        .O(\Q[26]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'hCCF0CC88FFFFFFFF)) 
    \Q[26]_i_14 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[28]_i_18_n_0 ),
        .I2(\Q[35]_i_20_n_0 ),
        .I3(\Q[17]_i_14_n_0 ),
        .I4(\Q[17]_i_11__0_n_0 ),
        .I5(\Q[22]_i_7__0_n_0 ),
        .O(\Q[26]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[26]_i_14__0 
       (.I0(\Q[35]_i_26_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[26]_i_14__0_n_0 ));
  LUT5 #(
    .INIT(32'h30353F35)) 
    \Q[26]_i_15 
       (.I0(\Q[35]_i_21_n_0 ),
        .I1(\Q[35]_i_20_n_0 ),
        .I2(\Q[29]_i_10_n_0 ),
        .I3(\Q[28]_i_20_n_0 ),
        .I4(\Q[35]_i_19_n_0 ),
        .O(\Q[26]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \Q[26]_i_15__0 
       (.I0(\Q[35]_i_18_n_0 ),
        .I1(EX_RF_RD1[28]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[154]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\custom_alu/int2fp/INT_VAL0 [28]),
        .O(\Q[26]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h0101050100000501)) 
    \Q[26]_i_16 
       (.I0(INT0_carry_i_6_n_0),
        .I1(ALU_DIN1[24]),
        .I2(INT0_carry__3_i_6_n_0),
        .I3(ALU_DIN1[21]),
        .I4(ALU_DIN1[23]),
        .I5(ALU_DIN1[22]),
        .O(\Q[26]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF088)) 
    \Q[26]_i_16__0 
       (.I0(\Q[17]_i_14_n_0 ),
        .I1(\Q[29]_i_18__0_n_0 ),
        .I2(\Q[17]_i_15_n_0 ),
        .I3(\Q[17]_i_10__0_n_0 ),
        .I4(\Q[69]_i_16_n_0 ),
        .I5(\Q[28]_i_11_n_0 ),
        .O(\Q[26]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[26]_i_17 
       (.I0(ALU_DIN1[0]),
        .I1(\Q[35]_i_20_n_0 ),
        .I2(\Q[28]_i_18_n_0 ),
        .I3(\Q[47]_i_9_n_0 ),
        .I4(\Q[17]_i_11__0_n_0 ),
        .I5(\Q[35]_i_32_n_0 ),
        .O(\Q[26]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h303F3737)) 
    \Q[26]_i_17__0 
       (.I0(\Q[31]_i_11__0_n_0 ),
        .I1(\Q[31]_i_13__0_n_0 ),
        .I2(\Q[29]_i_10_n_0 ),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[28]_i_20_n_0 ),
        .O(\Q[26]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h5555555533300030)) 
    \Q[26]_i_18 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_28_n_0 ),
        .I2(ALU_DIN1[17]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [17]),
        .I5(\Q[28]_i_11_n_0 ),
        .O(\Q[26]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h3353335F)) 
    \Q[26]_i_18__0 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[69]_i_16_n_0 ),
        .O(\Q[26]_i_18__0_n_0 ));
  LUT5 #(
    .INIT(32'hEFEC2020)) 
    \Q[26]_i_19 
       (.I0(\Q[29]_i_10_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[28]_i_20_n_0 ),
        .I4(\Q[23]_i_13__0_n_0 ),
        .O(\Q[26]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA6AAAAAA)) 
    \Q[26]_i_1__0 
       (.I0(\custom_alu/fp32_add/p_0_in [2]),
        .I1(\custom_alu/fp32_add/p_0_in [0]),
        .I2(\Q[30]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/significand_add0 [24]),
        .I4(\custom_alu/fp32_add/p_0_in [1]),
        .O(\custom_alu/fp32_add/p_1_out [26]));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[26]_i_1__1 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[27] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [3]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [26]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[26]_i_1__2 
       (.I0(\Q[26]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[11]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[11]),
        .I5(\Q[26]_i_4__0_n_0 ),
        .O(ID_RD2_FORWARDED[11]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[26]_i_1__3 
       (.I0(\Q[26]_i_2_n_0 ),
        .I1(\Q[26]_i_3__0_n_0 ),
        .I2(\Q[26]_i_4_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[21]),
        .O(data0[21]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[26]_i_1__4 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[26]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[21]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[26]_i_1__5 
       (.I0(ID_EX_Q[105]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[26]),
        .O(ALU_DIN2[26]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[26]_i_2 
       (.I0(\custom_alu/MULT [21]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [53]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [21]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEFEFFFFAEFEA)) 
    \Q[26]_i_20 
       (.I0(\Q[17]_i_14_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [13]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN1[13]),
        .I4(\custom_alu/int2fp/INT_VAL0 [14]),
        .I5(ALU_DIN1[14]),
        .O(\Q[26]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFAC00AF)) 
    \Q[26]_i_21 
       (.I0(\Q[29]_i_18__0_n_0 ),
        .I1(\Q[35]_i_32_n_0 ),
        .I2(\Q[35]_i_28_n_0 ),
        .I3(\Q[35]_i_29_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .O(\Q[26]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \Q[26]_i_22 
       (.I0(\Q[17]_i_15_n_0 ),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[35]_i_28_n_0 ),
        .I3(\Q[29]_i_18__0_n_0 ),
        .I4(\Q[47]_i_9_n_0 ),
        .O(\Q[26]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000511110005)) 
    \Q[26]_i_23 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [11]),
        .I2(ALU_DIN1[11]),
        .I3(ALU_DIN1[10]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [10]),
        .O(\Q[26]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[26]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[11]),
        .I2(CRF_RD2_IBUF[11]),
        .I3(RF_RD2_IBUF[11]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[26]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAFBAAAAAAAA)) 
    \Q[26]_i_3 
       (.I0(\Q[16]_i_2__0_n_0 ),
        .I1(\Q[26]_i_5__0_n_0 ),
        .I2(\Q[26]_i_6_n_0 ),
        .I3(EX_CUSTOM_ALU_SEL[28]),
        .I4(\Q[26]_i_7__0_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[11]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \Q[26]_i_3__0 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [21]),
        .O(\Q[26]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF8A88)) 
    \Q[26]_i_4 
       (.I0(EX_CUSTOM_ALU_SEL[26]),
        .I1(\Q[26]_i_5_n_0 ),
        .I2(\Q[26]_i_6__0_n_0 ),
        .I3(\Q[26]_i_7_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\Q[26]_i_8__0_n_0 ),
        .O(\Q[26]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \Q[26]_i_4__0 
       (.I0(DIN2_FORWARD[0]),
        .I1(DIN2_FORWARD[1]),
        .I2(data1[11]),
        .O(\Q[26]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFCA00C0)) 
    \Q[26]_i_5 
       (.I0(\Q[28]_i_12_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[28]_i_6_n_0 ),
        .I4(\Q[35]_i_16_n_0 ),
        .O(\Q[26]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEFEAFFFF)) 
    \Q[26]_i_5__0 
       (.I0(\custom_alu/fp2int/p_0_in [11]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I3(EX_RF_RD1[31]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[26]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA20000)) 
    \Q[26]_i_6 
       (.I0(\Q[26]_i_7_n_0 ),
        .I1(\Q[26]_i_9_n_0 ),
        .I2(\Q[26]_i_10__0_n_0 ),
        .I3(\Q[26]_i_11__0_n_0 ),
        .I4(\Q[27]_i_7_n_0 ),
        .I5(\Q[16]_i_4__1_n_0 ),
        .O(\Q[26]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88888888A8A8A8AA)) 
    \Q[26]_i_6__0 
       (.I0(\Q[26]_i_9__0_n_0 ),
        .I1(\Q[26]_i_10_n_0 ),
        .I2(\Q[26]_i_11_n_0 ),
        .I3(\Q[26]_i_12__0_n_0 ),
        .I4(\Q[26]_i_13__0_n_0 ),
        .I5(\Q[26]_i_14_n_0 ),
        .O(\Q[26]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000001DFF1D)) 
    \Q[26]_i_7 
       (.I0(EX_RF_RD1[30]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[156]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [30]),
        .I5(\Q[26]_i_15__0_n_0 ),
        .O(\Q[26]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \Q[26]_i_7__0 
       (.I0(\Q[69]_i_13_n_0 ),
        .I1(\Q[69]_i_14_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\custom_alu/fp32_mult/product_mantissa [11]),
        .I4(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .O(\Q[26]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    \Q[26]_i_8 
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__1_i_6_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__1_i_7_n_0),
        .O(\custom_alu/fp2int/p_0_in [11]));
  LUT5 #(
    .INIT(32'hFFFF3050)) 
    \Q[26]_i_8__0 
       (.I0(\Q[26]_i_16_n_0 ),
        .I1(\custom_alu/fp2int/INT0 [21]),
        .I2(EX_CUSTOM_ALU_SEL[27]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(EX_CUSTOM_ALU_SEL[28]),
        .O(\Q[26]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBABABABBBA)) 
    \Q[26]_i_9 
       (.I0(\Q[26]_i_12_n_0 ),
        .I1(\Q[26]_i_13_n_0 ),
        .I2(\Q[29]_i_7_n_0 ),
        .I3(\Q[26]_i_14__0_n_0 ),
        .I4(\Q[67]_i_12_n_0 ),
        .I5(\Q[26]_i_15_n_0 ),
        .O(\Q[26]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFA8)) 
    \Q[26]_i_9__0 
       (.I0(\Q[26]_i_17__0_n_0 ),
        .I1(\Q[26]_i_18__0_n_0 ),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[29]_i_7_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[26]_i_19_n_0 ),
        .O(\Q[26]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[27]_i_1 
       (.I0(\Q[27]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[28]),
        .O(CUSTOM_ALU_SEL[27]));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \Q[27]_i_13 
       (.I0(\Q[28]_i_20_n_0 ),
        .I1(\Q[28]_i_13_n_0 ),
        .I2(\Q[29]_i_7_n_0 ),
        .I3(\Q[35]_i_17_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[29]_i_13__0_n_0 ),
        .O(\Q[27]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h35373436FFFFFFFF)) 
    \Q[27]_i_14 
       (.I0(\Q[35]_i_26_n_0 ),
        .I1(\Q[35]_i_27_n_0 ),
        .I2(\Q[35]_i_22_n_0 ),
        .I3(\Q[35]_i_29_n_0 ),
        .I4(\Q[69]_i_21_n_0 ),
        .I5(\Q[69]_i_20_n_0 ),
        .O(\Q[27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF0F00FFFF22)) 
    \Q[27]_i_15 
       (.I0(\Q[69]_i_19_n_0 ),
        .I1(\Q[69]_i_18_n_0 ),
        .I2(\Q[17]_i_14_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[69]_i_16_n_0 ),
        .I5(\Q[17]_i_10__0_n_0 ),
        .O(\Q[27]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[27]_i_16 
       (.I0(exponent_carry_i_9_n_4),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_9_n_5),
        .O(\Q[27]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[27]_i_17 
       (.I0(exponent_carry_i_9_n_5),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_9_n_6),
        .O(\Q[27]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[27]_i_18 
       (.I0(exponent_carry_i_9_n_6),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_9_n_7),
        .O(\Q[27]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAA6AAAAAAAAAAAAA)) 
    \Q[27]_i_1__0 
       (.I0(\custom_alu/fp32_add/p_0_in [3]),
        .I1(\custom_alu/fp32_add/p_0_in [1]),
        .I2(\custom_alu/fp32_add/significand_add0 [24]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .I4(\custom_alu/fp32_add/p_0_in [0]),
        .I5(\custom_alu/fp32_add/p_0_in [2]),
        .O(\custom_alu/fp32_add/p_1_out [27]));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[27]_i_1__1 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[28] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [4]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [27]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[27]_i_1__2 
       (.I0(\Q[27]_i_2__1_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[12]),
        .I3(data1[12]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[12]));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[27]_i_1__3 
       (.I0(\Q[27]_i_2__0_n_0 ),
        .I1(\Q[27]_i_3__0_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[22]),
        .O(data0[22]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[27]_i_1__4 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[27]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[22]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[27]_i_1__5 
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[27]),
        .O(ALU_DIN2[27]));
  LUT5 #(
    .INIT(32'h10000000)) 
    \Q[27]_i_2 
       (.I0(CRF_RA2_OBUF[0]),
        .I1(CRF_RA2_OBUF[1]),
        .I2(\Q[29]_i_3_n_0 ),
        .I3(I_MEM_DOUT_IBUF[31]),
        .I4(\Q[27]_i_3_n_0 ),
        .O(\Q[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[27]_i_2__0 
       (.I0(\custom_alu/MULT [22]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [54]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(\custom_alu/Q [22]),
        .O(\Q[27]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[27]_i_2__1 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[12]),
        .I2(CRF_RD2_IBUF[12]),
        .I3(RF_RD2_IBUF[12]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[27]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \Q[27]_i_3 
       (.I0(CRF_RA2_OBUF[4]),
        .I1(I_MEM_DOUT_IBUF[30]),
        .I2(CRF_RA2_OBUF[3]),
        .I3(CRF_RA2_OBUF[2]),
        .O(\Q[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A0000FF8AFF8A)) 
    \Q[27]_i_3__0 
       (.I0(\Q[69]_i_5_n_0 ),
        .I1(\Q[27]_i_6_n_0 ),
        .I2(\Q[27]_i_7_n_0 ),
        .I3(EX_CUSTOM_ALU_SEL[28]),
        .I4(\Q[65]_i_5_n_0 ),
        .I5(\custom_alu/fp32_mult/product_mantissa [22]),
        .O(\Q[27]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h2A2A2A222A222A22)) 
    \Q[27]_i_6 
       (.I0(\Q[69]_i_12_n_0 ),
        .I1(\Q[26]_i_7_n_0 ),
        .I2(\Q[69]_i_11_n_0 ),
        .I3(\Q[27]_i_13_n_0 ),
        .I4(\Q[27]_i_14_n_0 ),
        .I5(\Q[27]_i_15_n_0 ),
        .O(\Q[27]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[27]_i_7 
       (.I0(EX_CUSTOM_ALU_SEL[26]),
        .I1(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[27]_i_7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[28]_i_1 
       (.I0(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .I1(I_MEM_DOUT_IBUF[28]),
        .O(CUSTOM_ALU_SEL[28]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF04)) 
    \Q[28]_i_10 
       (.I0(\Q[29]_i_10_n_0 ),
        .I1(\Q[28]_i_20_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[28]_i_21_n_0 ),
        .I4(\Q[35]_i_18_n_0 ),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[28]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[28]_i_11 
       (.I0(\custom_alu/int2fp/INT_VAL0 [18]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[144]),
        .I5(EX_RF_RD1[18]),
        .O(\Q[28]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[28]_i_12 
       (.I0(\custom_alu/int2fp/INT_VAL0 [26]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[152]),
        .I5(EX_RF_RD1[26]),
        .O(\Q[28]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \Q[28]_i_13 
       (.I0(ALU_DIN1[24]),
        .I1(\custom_alu/int2fp/INT_VAL0 [24]),
        .I2(ALU_DIN1[22]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [22]),
        .O(\Q[28]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \Q[28]_i_14 
       (.I0(\Q[17]_i_10__0_n_0 ),
        .I1(\Q[17]_i_14_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[31]_i_10__0_n_0 ),
        .O(\Q[28]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEAEAAFAAEFEA)) 
    \Q[28]_i_15 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [10]),
        .I2(\Q[63]_i_1__1_n_0 ),
        .I3(ALU_DIN1[10]),
        .I4(\custom_alu/int2fp/INT_VAL0 [11]),
        .I5(ALU_DIN1[11]),
        .O(\Q[28]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000001DFF1D)) 
    \Q[28]_i_16 
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[137]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [11]),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[28]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF4044)) 
    \Q[28]_i_17 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[28]_i_22_n_0 ),
        .I2(\Q[28]_i_23_n_0 ),
        .I3(\Q[28]_i_24_n_0 ),
        .I4(\Q[35]_i_26_n_0 ),
        .I5(\Q[35]_i_27_n_0 ),
        .O(\Q[28]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[28]_i_18 
       (.I0(\custom_alu/int2fp/INT_VAL0 [13]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[139]),
        .I5(EX_RF_RD1[13]),
        .O(\Q[28]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000001DFF1D)) 
    \Q[28]_i_19 
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [16]),
        .I5(\Q[17]_i_11__0_n_0 ),
        .O(\Q[28]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \Q[28]_i_1__0 
       (.I0(ALU_DIN1[27]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[27]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[106]),
        .I5(\Q[29]_i_2__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [28]));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[28]_i_1__1 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[29] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [5]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [28]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[28]_i_1__2 
       (.I0(\Q[28]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[13]),
        .I3(data1[13]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[13]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[28]_i_1__3 
       (.I0(\Q[28]_i_2_n_0 ),
        .I1(\Q[28]_i_3_n_0 ),
        .I2(\Q[28]_i_4_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[23]),
        .O(data0[23]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[28]_i_1__4 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[28]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[23]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[28]_i_1__5 
       (.I0(ID_EX_Q[107]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[28]),
        .O(ALU_DIN2[28]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[28]_i_2 
       (.I0(\custom_alu/MULT [23]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [55]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [23]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[28]_i_20 
       (.I0(\custom_alu/int2fp/INT_VAL0 [23]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[149]),
        .I5(EX_RF_RD1[23]),
        .O(\Q[28]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h000ACC0A)) 
    \Q[28]_i_21 
       (.I0(ALU_DIN1[25]),
        .I1(\custom_alu/int2fp/INT_VAL0 [25]),
        .I2(ALU_DIN1[26]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [26]),
        .O(\Q[28]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hCCAFFFAF)) 
    \Q[28]_i_22 
       (.I0(ALU_DIN1[5]),
        .I1(\custom_alu/int2fp/INT_VAL0 [5]),
        .I2(ALU_DIN1[4]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [4]),
        .O(\Q[28]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \Q[28]_i_23 
       (.I0(ALU_DIN1[5]),
        .I1(\custom_alu/int2fp/INT_VAL0 [5]),
        .I2(ALU_DIN1[3]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [3]),
        .O(\Q[28]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hCFAACFFFCCAACCAA)) 
    \Q[28]_i_24 
       (.I0(ALU_DIN1[2]),
        .I1(\custom_alu/int2fp/INT_VAL0 [2]),
        .I2(\custom_alu/int2fp/INT_VAL0 [1]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN1[1]),
        .I5(ALU_DIN1[0]),
        .O(\Q[28]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[28]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[13]),
        .I2(CRF_RD2_IBUF[13]),
        .I3(RF_RD2_IBUF[13]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[28]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[28]_i_2__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[28]),
        .I2(STALL_EN),
        .I3(IF_PC2[28]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[28] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[28]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h1F1F1F00)) 
    \Q[28]_i_3 
       (.I0(\custom_alu/fp32_mult/exponent_carry_n_7 ),
        .I1(\Q[35]_i_10_n_0 ),
        .I2(\Q[35]_i_11_n_0 ),
        .I3(\Q[28]_i_5_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[28]),
        .O(\Q[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[28]_i_3__0 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[27]),
        .I2(STALL_EN),
        .I3(IF_PC2[27]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[27] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[28]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8AAA8AAAA)) 
    \Q[28]_i_4 
       (.I0(\Q[30]_i_5_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[28]_i_7_n_0 ),
        .I3(\Q[28]_i_8_n_0 ),
        .I4(\Q[28]_i_9_n_0 ),
        .I5(\Q[28]_i_10_n_0 ),
        .O(\Q[28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[28]_i_4__0 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[26]),
        .I2(STALL_EN),
        .I3(IF_PC2[26]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[26] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[28]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h00FDFFFFFFFDFFFF)) 
    \Q[28]_i_5 
       (.I0(ALU_DIN1[24]),
        .I1(ALU_DIN1[23]),
        .I2(INT0_carry__4_i_4_n_0),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [23]),
        .O(\Q[28]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[28]_i_5__0 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[25]),
        .I2(STALL_EN),
        .I3(IF_PC2[25]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[25] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[28]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[28]_i_6 
       (.I0(\custom_alu/int2fp/INT_VAL0 [30]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[156]),
        .I5(EX_RF_RD1[30]),
        .O(\Q[28]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h000ACC0A)) 
    \Q[28]_i_7 
       (.I0(ALU_DIN1[28]),
        .I1(\custom_alu/int2fp/INT_VAL0 [28]),
        .I2(ALU_DIN1[29]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [29]),
        .O(\Q[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0F0FFF4)) 
    \Q[28]_i_8 
       (.I0(\Q[31]_i_10__0_n_0 ),
        .I1(\Q[28]_i_11_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[31]_i_11__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[28]_i_13_n_0 ),
        .O(\Q[28]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBBABAAAAAAAA)) 
    \Q[28]_i_9 
       (.I0(\Q[28]_i_14_n_0 ),
        .I1(\Q[28]_i_15_n_0 ),
        .I2(\Q[28]_i_16_n_0 ),
        .I3(\Q[28]_i_17_n_0 ),
        .I4(\Q[28]_i_18_n_0 ),
        .I5(\Q[28]_i_19_n_0 ),
        .O(\Q[28]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[29]_i_1 
       (.I0(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .I1(I_MEM_DOUT_IBUF[28]),
        .O(CUSTOM_ALU_SEL[29]));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[29]_i_10 
       (.I0(\custom_alu/int2fp/INT_VAL0 [24]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[150]),
        .I5(EX_RF_RD1[24]),
        .O(\Q[29]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h55544454FFFFFFFF)) 
    \Q[29]_i_10__0 
       (.I0(\Q[29]_i_16__0_n_0 ),
        .I1(\Q[66]_i_13_n_0 ),
        .I2(\Q[29]_i_17__0_n_0 ),
        .I3(\Q[35]_i_20_n_0 ),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[22]_i_7__0_n_0 ),
        .O(\Q[29]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT5 #(
    .INIT(32'hFFFFFF70)) 
    \Q[29]_i_11 
       (.I0(\Q[35]_i_22_n_0 ),
        .I1(ALU_DIN1[0]),
        .I2(\Q[69]_i_20_n_0 ),
        .I3(\Q[29]_i_19_n_0 ),
        .I4(\Q[27]_i_13_n_0 ),
        .O(\Q[29]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000001DFF1D)) 
    \Q[29]_i_11__0 
       (.I0(EX_RF_RD1[22]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[148]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [22]),
        .I5(\Q[31]_i_14__0_n_0 ),
        .O(\Q[29]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \Q[29]_i_12 
       (.I0(EX_RF_RD1[18]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[144]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [18]),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[29]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h5555555555554044)) 
    \Q[29]_i_12__0 
       (.I0(\Q[29]_i_19__0_n_0 ),
        .I1(\Q[29]_i_20_n_0 ),
        .I2(\Q[29]_i_21_n_0 ),
        .I3(\Q[29]_i_22_n_0 ),
        .I4(\Q[35]_i_21_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[29]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8B8B88B888888)) 
    \Q[29]_i_13 
       (.I0(\Q[17]_i_14_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[28]_i_18_n_0 ),
        .I4(\Q[31]_i_13__0_n_0 ),
        .I5(\Q[17]_i_11__0_n_0 ),
        .O(\Q[29]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00053305)) 
    \Q[29]_i_13__0 
       (.I0(ALU_DIN1[19]),
        .I1(\custom_alu/int2fp/INT_VAL0 [19]),
        .I2(ALU_DIN1[20]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [20]),
        .O(\Q[29]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000F77FFFF0F77)) 
    \Q[29]_i_14 
       (.I0(\Q[35]_i_21_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[35]_i_19_n_0 ),
        .I3(\Q[31]_i_11__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[35]_i_20_n_0 ),
        .O(\Q[29]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_15 
       (.I0(EX_RF_RD1[24]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[150]),
        .O(\Q[29]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \Q[29]_i_15__0 
       (.I0(\Q[17]_i_10__0_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[69]_i_16_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[29]_i_15__0_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_16 
       (.I0(EX_RF_RD1[23]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[149]),
        .O(\Q[29]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h5555303F55553030)) 
    \Q[29]_i_16__0 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_28_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[17]_i_15_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[29]_i_16__0_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_17 
       (.I0(EX_RF_RD1[22]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[148]),
        .O(\custom_alu/int2fp/INT_VAL1 [22]));
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \Q[29]_i_17__0 
       (.I0(\Q[35]_i_32_n_0 ),
        .I1(\Q[35]_i_19_n_0 ),
        .I2(ALU_DIN1[1]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [1]),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[29]_i_17__0_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_18 
       (.I0(EX_RF_RD1[21]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[147]),
        .O(\custom_alu/int2fp/INT_VAL1 [21]));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[29]_i_18__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [3]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[129]),
        .I5(EX_RF_RD1[3]),
        .O(\Q[29]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'h303F3535303F3030)) 
    \Q[29]_i_19 
       (.I0(\Q[35]_i_26_n_0 ),
        .I1(\Q[35]_i_22_n_0 ),
        .I2(\Q[28]_i_11_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[69]_i_16_n_0 ),
        .I5(\Q[17]_i_10__0_n_0 ),
        .O(\Q[29]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \Q[29]_i_19__0 
       (.I0(ALU_DIN1[11]),
        .I1(\custom_alu/int2fp/INT_VAL0 [11]),
        .I2(ALU_DIN1[12]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [12]),
        .O(\Q[29]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h3CCC5A5A3CCCAAAA)) 
    \Q[29]_i_1__0 
       (.I0(ALU_DIN1[28]),
        .I1(ALU_DIN2[28]),
        .I2(\Q[29]_i_2__0_n_0 ),
        .I3(ALU_DIN2[27]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN1[27]),
        .O(\custom_alu/fp32_add/p_1_out [29]));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[29]_i_1__1 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[30] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [6]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [29]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[29]_i_1__2 
       (.I0(\Q[29]_i_2__2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[14]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[14]),
        .I5(\Q[29]_i_4__1_n_0 ),
        .O(ID_RD2_FORWARDED[14]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[29]_i_1__3 
       (.I0(\Q[29]_i_2__1_n_0 ),
        .I1(\Q[29]_i_3__1_n_0 ),
        .I2(\Q[29]_i_4__0_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[24]),
        .O(data0[24]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[29]_i_1__4 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[29]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[24]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[24]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[29]_i_1__5 
       (.I0(ID_EX_Q[108]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[29]),
        .O(ALU_DIN2[29]));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \Q[29]_i_2 
       (.I0(I_MEM_DOUT_IBUF[31]),
        .I1(I_MEM_DOUT_IBUF[30]),
        .I2(\Q[29]_i_3_n_0 ),
        .O(CUSTOM_INSTRUCTION_STALL_CYCLE[1]));
  LUT5 #(
    .INIT(32'h00053305)) 
    \Q[29]_i_20 
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/int2fp/INT_VAL0 [7]),
        .I2(ALU_DIN1[8]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [8]),
        .O(\Q[29]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFE200E2)) 
    \Q[29]_i_21 
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [5]),
        .I5(\Q[35]_i_29_n_0 ),
        .O(\Q[29]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF04)) 
    \Q[29]_i_22 
       (.I0(\Q[35]_i_32_n_0 ),
        .I1(ALU_DIN1[0]),
        .I2(\Q[47]_i_9_n_0 ),
        .I3(\Q[29]_i_18__0_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .O(\Q[29]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_23 
       (.I0(EX_RF_RD1[28]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[154]),
        .O(\Q[29]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_24 
       (.I0(EX_RF_RD1[27]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[153]),
        .O(\Q[29]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_25 
       (.I0(EX_RF_RD1[26]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[152]),
        .O(\Q[29]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[29]_i_26 
       (.I0(EX_RF_RD1[25]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[151]),
        .O(\Q[29]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \Q[29]_i_2__0 
       (.I0(\custom_alu/fp32_add/p_0_in [3]),
        .I1(\custom_alu/fp32_add/p_0_in [1]),
        .I2(\custom_alu/fp32_add/significand_add0 [24]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .I4(\custom_alu/fp32_add/p_0_in [0]),
        .I5(\custom_alu/fp32_add/p_0_in [2]),
        .O(\Q[29]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[29]_i_2__1 
       (.I0(\custom_alu/MULT [24]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [56]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [24]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[29]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[29]_i_2__2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[14]),
        .I2(CRF_RD2_IBUF[14]),
        .I3(RF_RD2_IBUF[14]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[29]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    \Q[29]_i_3 
       (.I0(I_MEM_DOUT_IBUF[6]),
        .I1(I_MEM_DOUT_IBUF[3]),
        .I2(\Q[29]_i_4_n_0 ),
        .I3(I_MEM_DOUT_IBUF[25]),
        .I4(EX_BR_TAKEN),
        .I5(I_MEM_DOUT_IBUF[5]),
        .O(\Q[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF10FFFFFF100000)) 
    \Q[29]_i_3__0 
       (.I0(\Q[29]_i_5_n_0 ),
        .I1(\Q[29]_i_6__0_n_0 ),
        .I2(\Q[29]_i_7__0_n_0 ),
        .I3(\Q[29]_i_8__0_n_0 ),
        .I4(\Q[34]_i_5_n_0 ),
        .I5(\Q[19]_i_3__0_n_0 ),
        .O(CUSTOM_ALU_OUT[14]));
  LUT6 #(
    .INIT(64'hF200FFFFFFFFFFFF)) 
    \Q[29]_i_3__1 
       (.I0(\Q[29]_i_5__0_n_0 ),
        .I1(\Q[29]_i_6_n_0 ),
        .I2(\Q[29]_i_7_n_0 ),
        .I3(\Q[29]_i_8_n_0 ),
        .I4(\Q[30]_i_5__0_n_0 ),
        .I5(\Q[30]_i_5_n_0 ),
        .O(\Q[29]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000005510)) 
    \Q[29]_i_4 
       (.I0(I_MEM_DOUT_IBUF[29]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(I_MEM_DOUT_IBUF[4]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[27]),
        .I5(I_MEM_DOUT_IBUF[26]),
        .O(\Q[29]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT4 #(
    .INIT(16'hFEAA)) 
    \Q[29]_i_4__0 
       (.I0(\Q[30]_i_2__0_n_0 ),
        .I1(\custom_alu/fp32_mult/exponent_carry_n_6 ),
        .I2(\Q[35]_i_10_n_0 ),
        .I3(\Q[35]_i_11_n_0 ),
        .O(\Q[29]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \Q[29]_i_4__1 
       (.I0(DIN2_FORWARD[0]),
        .I1(DIN2_FORWARD[1]),
        .I2(data1[14]),
        .O(\Q[29]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555DD5D)) 
    \Q[29]_i_5 
       (.I0(\Q[26]_i_7_n_0 ),
        .I1(\Q[29]_i_9_n_0 ),
        .I2(\Q[29]_i_10__0_n_0 ),
        .I3(\Q[29]_i_11_n_0 ),
        .I4(\Q[29]_i_12_n_0 ),
        .I5(\Q[19]_i_4__0_n_0 ),
        .O(\Q[29]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000001DFF1D)) 
    \Q[29]_i_5__0 
       (.I0(EX_RF_RD1[23]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[149]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [23]),
        .I5(\Q[29]_i_10_n_0 ),
        .O(\Q[29]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880008AAAAAAAA)) 
    \Q[29]_i_6 
       (.I0(\Q[29]_i_11__0_n_0 ),
        .I1(\Q[31]_i_12__0_n_0 ),
        .I2(\Q[35]_i_24_n_0 ),
        .I3(\Q[29]_i_12__0_n_0 ),
        .I4(\Q[35]_i_23_n_0 ),
        .I5(\Q[29]_i_13__0_n_0 ),
        .O(\Q[29]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[29]_i_6__0 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [14]),
        .O(\Q[29]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \Q[29]_i_7 
       (.I0(ALU_DIN1[25]),
        .I1(\custom_alu/int2fp/INT_VAL0 [25]),
        .I2(ALU_DIN1[26]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [26]),
        .O(\Q[29]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hEFEAFFFF)) 
    \Q[29]_i_7__0 
       (.I0(INT0_carry__2_i_8_n_0),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[29]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000015155550151)) 
    \Q[29]_i_8 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(EX_RF_RD1[28]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[154]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [28]),
        .O(\Q[29]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \Q[29]_i_8__0 
       (.I0(\Q[69]_i_13_n_0 ),
        .I1(\Q[69]_i_14_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\custom_alu/fp32_mult/product_mantissa [14]),
        .I4(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .O(\Q[29]_i_8__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1110)) 
    \Q[29]_i_9 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[29]_i_13_n_0 ),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[29]_i_14_n_0 ),
        .I4(\Q[29]_i_15__0_n_0 ),
        .O(\Q[29]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[2]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [1]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [2]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [2]));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[2]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[3] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/data23 [2]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\Q[2]_i_2_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [2]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[2]_i_1__1 
       (.I0(I_MEM_DOUT_IBUF[9]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[9]));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT4 #(
    .INIT(16'h0708)) 
    \Q[2]_i_1__2 
       (.I0(STALL_COUNTER_Q[1]),
        .I1(STALL_COUNTER_Q[0]),
        .I2(STALL_COUNTER_D1),
        .I3(STALL_COUNTER_Q[2]),
        .O(STALL_COUNTER_D[2]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[2]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [0]),
        .O(\Q[2]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT4 #(
    .INIT(16'h0200)) 
    \Q[30]_i_1 
       (.I0(\Q[31]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[14]),
        .I2(I_MEM_DOUT_IBUF[13]),
        .I3(I_MEM_DOUT_IBUF[12]),
        .O(CUSTOM_ALU_SEL[30]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4700)) 
    \Q[30]_i_10 
       (.I0(\Q[47]_i_9_n_0 ),
        .I1(\Q[35]_i_22_n_0 ),
        .I2(\Q[30]_i_17_n_0 ),
        .I3(\Q[69]_i_20_n_0 ),
        .I4(\Q[20]_i_13__0_n_0 ),
        .I5(\Q[27]_i_13_n_0 ),
        .O(\Q[30]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000110111111111)) 
    \Q[30]_i_10__0 
       (.I0(\Q[35]_i_23_n_0 ),
        .I1(\Q[35]_i_24_n_0 ),
        .I2(ALU_DIN1[0]),
        .I3(\Q[35]_i_25_n_0 ),
        .I4(\Q[30]_i_13__0_n_0 ),
        .I5(\Q[30]_i_14_n_0 ),
        .O(\Q[30]_i_10__0_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[30]_i_11 
       (.I0(EX_RF_RD1[30]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[156]),
        .O(\Q[30]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \Q[30]_i_11__0 
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[145]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [19]),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[30]_i_11__0_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[30]_i_12 
       (.I0(EX_RF_RD1[29]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[155]),
        .O(\Q[30]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8B8B88B888888)) 
    \Q[30]_i_12__0 
       (.I0(\Q[17]_i_10__0_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[17]_i_11__0_n_0 ),
        .I4(\Q[31]_i_13__0_n_0 ),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[30]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000F77FFFF0F77)) 
    \Q[30]_i_13 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[35]_i_20_n_0 ),
        .I3(\Q[31]_i_11__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[30]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFEFEFE)) 
    \Q[30]_i_13__0 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_28_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\custom_alu/int2fp/INT_VAL0 [7]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN1[7]),
        .O(\Q[30]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001015)) 
    \Q[30]_i_14 
       (.I0(\Q[35]_i_22_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [10]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN1[10]),
        .I4(\Q[35]_i_20_n_0 ),
        .I5(\Q[35]_i_19_n_0 ),
        .O(\Q[30]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \Q[30]_i_14__0 
       (.I0(\Q[69]_i_16_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[30]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'h5555303F55553030)) 
    \Q[30]_i_15 
       (.I0(\Q[35]_i_26_n_0 ),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[35]_i_28_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[30]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \Q[30]_i_16 
       (.I0(\Q[29]_i_18__0_n_0 ),
        .I1(\Q[35]_i_19_n_0 ),
        .I2(ALU_DIN1[2]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [2]),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[30]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \Q[30]_i_17 
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[134]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [8]),
        .I5(ALU_DIN1[0]),
        .O(\Q[30]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[30]_i_19 
       (.I0(EX_RF_RD1[20]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[146]),
        .O(\custom_alu/int2fp/INT_VAL1 [20]));
  LUT6 #(
    .INIT(64'hFFFF7FFF00008000)) 
    \Q[30]_i_1__0 
       (.I0(\custom_alu/fp32_add/p_0_in [4]),
        .I1(\Q[30]_i_2_n_0 ),
        .I2(\custom_alu/fp32_add/p_0_in [5]),
        .I3(\custom_alu/fp32_add/significand_add0 [24]),
        .I4(\Q[30]_i_4__0_n_0 ),
        .I5(\custom_alu/fp32_add/p_0_in [6]),
        .O(\custom_alu/fp32_add/p_1_out [30]));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[30]_i_1__1 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[31] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/exp_sub [7]),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [30]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[30]_i_1__2 
       (.I0(\Q[30]_i_2__2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[15]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[15]),
        .I5(\Q[30]_i_4__1_n_0 ),
        .O(ID_RD2_FORWARDED[15]));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \Q[30]_i_1__3 
       (.I0(\Q[30]_i_2__0_n_0 ),
        .I1(\Q[30]_i_3__0_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\Q[30]_i_4_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[25]),
        .O(data0[25]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[30]_i_1__4 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[30]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[25]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[25]));
  LUT2 #(
    .INIT(4'hB)) 
    \Q[30]_i_1__5 
       (.I0(IF_PC_ADD4[30]),
        .I1(RSTn_IBUF),
        .O(D0));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[30]_i_1__6 
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[30]),
        .O(ALU_DIN2[30]));
  LUT6 #(
    .INIT(64'hB800000000000000)) 
    \Q[30]_i_2 
       (.I0(ALU_DIN2[23]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[23]),
        .I3(\custom_alu/fp32_add/p_0_in [1]),
        .I4(\custom_alu/fp32_add/p_0_in [3]),
        .I5(\custom_alu/fp32_add/p_0_in [2]),
        .O(\Q[30]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[30]_i_20 
       (.I0(EX_RF_RD1[19]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[145]),
        .O(\custom_alu/int2fp/INT_VAL1 [19]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[30]_i_21 
       (.I0(EX_RF_RD1[18]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[144]),
        .O(\custom_alu/int2fp/INT_VAL1 [18]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[30]_i_22 
       (.I0(EX_RF_RD1[17]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[143]),
        .O(\Q[30]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000045400000)) 
    \Q[30]_i_2__0 
       (.I0(\custom_alu/fp2int/INT0_carry__4_n_0 ),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(EX_CUSTOM_ALU_SEL[28]),
        .O(\Q[30]_i_2__0_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2)) 
    \Q[30]_i_2__1 
       (.I0(EX_RF_RD2[31]),
        .I1(\FF_ID_EX/Q_reg_n_0_[158] ),
        .I2(ID_EX_Q[110]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .O(\Q[30]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[30]_i_2__2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[15]),
        .I2(CRF_RD2_IBUF[15]),
        .I3(RF_RD2_IBUF[15]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[30]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBBFBAAAAAAAA)) 
    \Q[30]_i_3 
       (.I0(\Q[20]_i_2__0_n_0 ),
        .I1(\Q[20]_i_3__1_n_0 ),
        .I2(\Q[30]_i_5_n_0 ),
        .I3(\Q[30]_i_6_n_0 ),
        .I4(\Q[30]_i_7_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[15]));
  LUT6 #(
    .INIT(64'hFFFFFFD0D0D0D0D0)) 
    \Q[30]_i_3__0 
       (.I0(\Q[30]_i_5__0_n_0 ),
        .I1(\Q[30]_i_6__0_n_0 ),
        .I2(\Q[30]_i_5_n_0 ),
        .I3(\custom_alu/fp32_mult/exponent_carry_n_5 ),
        .I4(\Q[35]_i_10_n_0 ),
        .I5(\Q[35]_i_11_n_0 ),
        .O(\Q[30]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[30]_i_4 
       (.I0(\custom_alu/MULT [25]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [57]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(\custom_alu/Q [25]),
        .O(\Q[30]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hBEBBBEEE)) 
    \Q[30]_i_4__0 
       (.I0(\Q[88]_i_3_n_0 ),
        .I1(PSUM3__0_carry__0_i_10__2_n_0),
        .I2(ID_EX_Q[110]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[31]),
        .O(\Q[30]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \Q[30]_i_4__1 
       (.I0(DIN2_FORWARD[0]),
        .I1(DIN2_FORWARD[1]),
        .I2(data1[15]),
        .O(\Q[30]_i_4__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \Q[30]_i_5 
       (.I0(EX_CUSTOM_ALU_SEL[27]),
        .I1(EX_CUSTOM_ALU_SEL[26]),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .O(\Q[30]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000015155550151)) 
    \Q[30]_i_5__0 
       (.I0(\Q[28]_i_6_n_0 ),
        .I1(EX_RF_RD1[29]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[155]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [29]),
        .O(\Q[30]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h00008808AAAAAAAA)) 
    \Q[30]_i_6 
       (.I0(\Q[20]_i_7__0_n_0 ),
        .I1(\Q[30]_i_8_n_0 ),
        .I2(\Q[30]_i_9__0_n_0 ),
        .I3(\Q[30]_i_10_n_0 ),
        .I4(\Q[30]_i_11__0_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[30]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAA08AA)) 
    \Q[30]_i_6__0 
       (.I0(\Q[30]_i_8__0_n_0 ),
        .I1(\Q[30]_i_9_n_0 ),
        .I2(\Q[30]_i_10__0_n_0 ),
        .I3(\Q[29]_i_5__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[31]_i_13__0_n_0 ),
        .O(\Q[30]_i_6__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \Q[30]_i_7 
       (.I0(\Q[69]_i_13_n_0 ),
        .I1(\Q[69]_i_14_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\custom_alu/fp32_mult/product_mantissa [15]),
        .I4(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .O(\Q[30]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1110)) 
    \Q[30]_i_8 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[30]_i_12__0_n_0 ),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[30]_i_13_n_0 ),
        .I4(\Q[30]_i_14__0_n_0 ),
        .O(\Q[30]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000047)) 
    \Q[30]_i_8__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [28]),
        .I1(PSUM3__0_carry__0_i_10__2_n_0),
        .I2(ALU_DIN1[28]),
        .I3(\Q[35]_i_17_n_0 ),
        .I4(\Q[29]_i_7_n_0 ),
        .O(\Q[30]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000010101)) 
    \Q[30]_i_9 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\custom_alu/int2fp/INT_VAL0 [19]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(ALU_DIN1[19]),
        .O(\Q[30]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h55544454FFFFFFFF)) 
    \Q[30]_i_9__0 
       (.I0(\Q[30]_i_15_n_0 ),
        .I1(\Q[66]_i_13_n_0 ),
        .I2(\Q[30]_i_16_n_0 ),
        .I3(\Q[35]_i_20_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .I5(\Q[22]_i_7__0_n_0 ),
        .O(\Q[30]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \Q[31]_i_1 
       (.I0(\Q[31]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[12]),
        .I3(I_MEM_DOUT_IBUF[14]),
        .O(CUSTOM_ALU_SEL[31]));
  LUT6 #(
    .INIT(64'hB8FFB800B800B800)) 
    \Q[31]_i_10 
       (.I0(\custom_alu/int2fp/INT_VAL0 [4]),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN1[4]),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[35]_i_21_n_0 ),
        .O(\Q[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[31]_i_10__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [19]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[145]),
        .I5(EX_RF_RD1[19]),
        .O(\Q[31]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[31]_i_11 
       (.I0(\Q[35]_i_32_n_0 ),
        .I1(\Q[35]_i_22_n_0 ),
        .I2(\Q[47]_i_9_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(ALU_DIN1[0]),
        .I5(\Q[35]_i_26_n_0 ),
        .O(\Q[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[31]_i_11__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [20]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[146]),
        .I5(EX_RF_RD1[20]),
        .O(\Q[31]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h30353F3530303F30)) 
    \Q[31]_i_12 
       (.I0(\Q[35]_i_22_n_0 ),
        .I1(\Q[35]_i_19_n_0 ),
        .I2(\Q[28]_i_11_n_0 ),
        .I3(\Q[69]_i_16_n_0 ),
        .I4(\Q[35]_i_21_n_0 ),
        .I5(\Q[17]_i_10__0_n_0 ),
        .O(\Q[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000001DFF1D)) 
    \Q[31]_i_12__0 
       (.I0(EX_RF_RD1[17]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(ID_EX_Q[143]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [17]),
        .I5(\Q[28]_i_11_n_0 ),
        .O(\Q[31]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000F77FFFF0F77)) 
    \Q[31]_i_13 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[28]_i_18_n_0 ),
        .I3(\Q[31]_i_11__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[17]_i_11__0_n_0 ),
        .O(\Q[31]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[31]_i_13__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [22]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[148]),
        .I5(EX_RF_RD1[22]),
        .O(\Q[31]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEEAFAAAAEEAF)) 
    \Q[31]_i_14 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[31]_i_15_n_0 ),
        .I3(\Q[28]_i_20_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[69]_i_16_n_0 ),
        .O(\Q[31]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[31]_i_14__0 
       (.I0(\custom_alu/int2fp/INT_VAL0 [21]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[147]),
        .I5(EX_RF_RD1[21]),
        .O(\Q[31]_i_14__0_n_0 ));
  LUT5 #(
    .INIT(32'h335FFF5F)) 
    \Q[31]_i_15 
       (.I0(ALU_DIN1[22]),
        .I1(\custom_alu/int2fp/INT_VAL0 [22]),
        .I2(ALU_DIN1[15]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [15]),
        .O(\Q[31]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1DE2E2E2E2E2E2E2)) 
    \Q[31]_i_1__0 
       (.I0(ALU_DIN1[30]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN2[30]),
        .I3(\custom_alu/fp32_add/p_0_in [5]),
        .I4(\custom_alu/fp32_add/p_0_in [6]),
        .I5(\Q[31]_i_2__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [31]));
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[31]_i_1__1 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[0] ),
        .I1(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [31]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[31]_i_1__2 
       (.I0(\Q[31]_i_2__3_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[16]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[16]),
        .I5(\Q[31]_i_4__1_n_0 ),
        .O(ID_RD2_FORWARDED[16]));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \Q[31]_i_1__3 
       (.I0(\Q[31]_i_2__2_n_0 ),
        .I1(\Q[31]_i_3__2_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\Q[31]_i_4__0_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[26]),
        .O(data0[26]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[31]_i_1__4 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[31]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[26]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[26]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[31]_i_1__5 
       (.I0(ID_EX_Q[110]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[31]),
        .O(ALU_DIN2[31]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \Q[31]_i_2 
       (.I0(\Q[31]_i_3_n_0 ),
        .I1(\Q[161]_i_2_n_0 ),
        .I2(I_MEM_DOUT_IBUF[29]),
        .I3(\Q[123]_i_3_n_0 ),
        .I4(I_MEM_DOUT_IBUF[27]),
        .I5(I_MEM_DOUT_IBUF[26]),
        .O(\Q[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \Q[31]_i_2__0 
       (.I0(ALU_DIN1[27]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[27]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(ID_EX_Q[106]),
        .I5(\Q[29]_i_2__0_n_0 ),
        .O(\Q[31]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF80000000)) 
    \Q[31]_i_2__1 
       (.I0(\custom_alu/fp32_add/p_0_in [6]),
        .I1(\custom_alu/fp32_add/p_0_in [7]),
        .I2(\custom_alu/fp32_add/p_0_in [4]),
        .I3(\custom_alu/fp32_add/p_0_in [5]),
        .I4(\Q[30]_i_2_n_0 ),
        .I5(\Q[31]_i_3__0_n_0 ),
        .O(\Q[31]_i_2__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hA8)) 
    \Q[31]_i_2__2 
       (.I0(\Q[35]_i_11_n_0 ),
        .I1(\Q[35]_i_10_n_0 ),
        .I2(\custom_alu/fp32_mult/exponent_carry_n_4 ),
        .O(\Q[31]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[31]_i_2__3 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[16]),
        .I2(CRF_RD2_IBUF[16]),
        .I3(RF_RD2_IBUF[16]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[31]_i_2__3_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[31]_i_2__4 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[31]),
        .I2(STALL_EN),
        .I3(IF_PC2[31]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[31] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[31]_i_2__4_n_0 ));
  LUT6 #(
    .INIT(64'h0100010001000000)) 
    \Q[31]_i_3 
       (.I0(I_MEM_DOUT_IBUF[28]),
        .I1(I_MEM_DOUT_IBUF[30]),
        .I2(I_MEM_DOUT_IBUF[31]),
        .I3(I_MEM_DOUT_IBUF[25]),
        .I4(EX_BR_TAKEN),
        .I5(I_MEM_DOUT_IBUF[5]),
        .O(\Q[31]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \Q[31]_i_3__0 
       (.I0(\Q[31]_i_4_n_0 ),
        .I1(\custom_alu/fp32_add/p_0_in2_in [1]),
        .I2(\custom_alu/fp32_add/p_0_in2_in [2]),
        .I3(\custom_alu/fp32_add/p_0_in2_in [5]),
        .I4(\custom_alu/fp32_add/p_0_in2_in [6]),
        .O(\Q[31]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFFFBAAAAAAAA)) 
    \Q[31]_i_3__1 
       (.I0(\Q[21]_i_2__0_n_0 ),
        .I1(\Q[21]_i_3__0_n_0 ),
        .I2(\Q[31]_i_5_n_0 ),
        .I3(\custom_alu/fp32_mult/product_mantissa [16]),
        .I4(\Q[65]_i_5_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[16]));
  LUT6 #(
    .INIT(64'hFFBFBBBBAAAAAAAA)) 
    \Q[31]_i_3__2 
       (.I0(\Q[30]_i_2__0_n_0 ),
        .I1(\Q[31]_i_5__0_n_0 ),
        .I2(\Q[35]_i_8_n_0 ),
        .I3(\Q[31]_i_6__0_n_0 ),
        .I4(\Q[31]_i_7__0_n_0 ),
        .I5(\Q[30]_i_5_n_0 ),
        .O(\Q[31]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FFE4FFE4FF)) 
    \Q[31]_i_3__3 
       (.I0(EX_BR_TAKEN),
        .I1(\FF_IF_ID_PCADD/Q_reg_n_0_[30] ),
        .I2(IF_PC2[30]),
        .I3(RSTn_IBUF),
        .I4(ID_PC[30]),
        .I5(STALL_EN),
        .O(\Q[31]_i_3__3_n_0 ));
  LUT6 #(
    .INIT(64'h8000808080000000)) 
    \Q[31]_i_4 
       (.I0(\custom_alu/fp32_add/p_0_in2_in [3]),
        .I1(\custom_alu/fp32_add/p_0_in2_in [0]),
        .I2(\custom_alu/fp32_add/p_0_in2_in [4]),
        .I3(ALU_DIN1[30]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[30]),
        .O(\Q[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[31]_i_4__0 
       (.I0(\custom_alu/MULT [26]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [58]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(EX_CUSTOM_ALU_SEL[29]),
        .I5(\custom_alu/Q [26]),
        .O(\Q[31]_i_4__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \Q[31]_i_4__1 
       (.I0(DIN2_FORWARD[0]),
        .I1(DIN2_FORWARD[1]),
        .I2(data1[16]),
        .O(\Q[31]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[31]_i_4__2 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[29]),
        .I2(STALL_EN),
        .I3(IF_PC2[29]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[29] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[31]_i_4__2_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \Q[31]_i_5 
       (.I0(\Q[30]_i_5_n_0 ),
        .I1(\Q[21]_i_7__0_n_0 ),
        .I2(\Q[31]_i_6_n_0 ),
        .I3(\Q[31]_i_7_n_0 ),
        .I4(\Q[31]_i_8_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[31]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \Q[31]_i_5__0 
       (.I0(\Q[35]_i_18_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[29]_i_7_n_0 ),
        .I3(\Q[35]_i_17_n_0 ),
        .I4(\Q[35]_i_16_n_0 ),
        .O(\Q[31]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h55544454FFFFFFFF)) 
    \Q[31]_i_6 
       (.I0(\Q[31]_i_9_n_0 ),
        .I1(\Q[66]_i_13_n_0 ),
        .I2(\Q[31]_i_10_n_0 ),
        .I3(\Q[35]_i_20_n_0 ),
        .I4(\Q[35]_i_28_n_0 ),
        .I5(\Q[22]_i_7__0_n_0 ),
        .O(\Q[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \Q[31]_i_6__0 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_28_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[35]_i_25_n_0 ),
        .I5(ALU_DIN1[0]),
        .O(\Q[31]_i_6__0_n_0 ));
  LUT4 #(
    .INIT(16'hFFF4)) 
    \Q[31]_i_7 
       (.I0(\Q[31]_i_11_n_0 ),
        .I1(\Q[69]_i_20_n_0 ),
        .I2(\Q[31]_i_12_n_0 ),
        .I3(\Q[27]_i_13_n_0 ),
        .O(\Q[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \Q[31]_i_7__0 
       (.I0(\Q[31]_i_10__0_n_0 ),
        .I1(\Q[31]_i_11__0_n_0 ),
        .I2(\Q[31]_i_12__0_n_0 ),
        .I3(\Q[31]_i_13__0_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[29]_i_5__0_n_0 ),
        .O(\Q[31]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h7070707077777770)) 
    \Q[31]_i_8 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(\Q[31]_i_11__0_n_0 ),
        .I2(\Q[21]_i_9__0_n_0 ),
        .I3(\Q[31]_i_13_n_0 ),
        .I4(\Q[67]_i_12_n_0 ),
        .I5(\Q[31]_i_14_n_0 ),
        .O(\Q[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5555303F55553030)) 
    \Q[31]_i_9 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[35]_i_26_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[35]_i_29_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[31]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[32]_i_1 
       (.I0(\Q[32]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[17]),
        .I3(data1[17]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[17]));
  LUT5 #(
    .INIT(32'h8AFF8A00)) 
    \Q[32]_i_1__0 
       (.I0(\Q[32]_i_2_n_0 ),
        .I1(\Q[32]_i_3_n_0 ),
        .I2(\Q[32]_i_4_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[27]),
        .O(data0[27]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[32]_i_1__1 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[32]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[27]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[27]));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \Q[32]_i_2 
       (.I0(\custom_alu/Q [27]),
        .I1(EX_CUSTOM_ALU_SEL[29]),
        .I2(EX_CUSTOM_ALU_SEL[30]),
        .I3(\custom_alu/MULT [59]),
        .I4(EX_CUSTOM_ALU_SEL[31]),
        .I5(\custom_alu/MULT [27]),
        .O(\Q[32]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[32]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[17]),
        .I2(CRF_RD2_IBUF[17]),
        .I3(RF_RD2_IBUF[17]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[32]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFDFDDDD)) 
    \Q[32]_i_3 
       (.I0(\Q[34]_i_5_n_0 ),
        .I1(\Q[30]_i_2__0_n_0 ),
        .I2(\Q[35]_i_7_n_0 ),
        .I3(\Q[34]_i_6_n_0 ),
        .I4(\Q[30]_i_5_n_0 ),
        .O(\Q[32]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'h1F)) 
    \Q[32]_i_4 
       (.I0(\Q[35]_i_10_n_0 ),
        .I1(\custom_alu/fp32_mult/exponent_carry__0_n_7 ),
        .I2(\Q[35]_i_11_n_0 ),
        .O(\Q[32]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[33]_i_1 
       (.I0(\Q[33]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[18]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[18]),
        .I5(\Q[33]_i_3__0_n_0 ),
        .O(ID_RD2_FORWARDED[18]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[33]_i_1__0 
       (.I0(\Q[33]_i_2_n_0 ),
        .I1(\Q[34]_i_3_n_0 ),
        .I2(\Q[33]_i_3_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[28]),
        .O(data0[28]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[33]_i_1__1 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[33]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[28]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[28]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[33]_i_2 
       (.I0(\custom_alu/MULT [28]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [60]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [28]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[33]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[33]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[18]),
        .I2(CRF_RD2_IBUF[18]),
        .I3(RF_RD2_IBUF[18]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[33]_i_2__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hA8)) 
    \Q[33]_i_3 
       (.I0(\Q[35]_i_11_n_0 ),
        .I1(\Q[35]_i_10_n_0 ),
        .I2(\custom_alu/fp32_mult/exponent_carry__0_n_6 ),
        .O(\Q[33]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA80AA8080)) 
    \Q[33]_i_3__0 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(\Q[36]_i_3__0_n_0 ),
        .I2(D_MEM_DOUT_IBUF[18]),
        .I3(MEM_D_MEM_ALU_FINAL1),
        .I4(EX_MEM_Q[23]),
        .I5(\Q[36]_i_2__1_n_0 ),
        .O(\Q[33]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[34]_i_1 
       (.I0(\Q[34]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[19]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[19]),
        .I5(\Q[34]_i_3__0_n_0 ),
        .O(ID_RD2_FORWARDED[19]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[34]_i_1__0 
       (.I0(\Q[34]_i_2_n_0 ),
        .I1(\Q[34]_i_3_n_0 ),
        .I2(\Q[34]_i_4_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[29]),
        .O(data0[29]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[34]_i_1__1 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[34]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[29]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[29]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[34]_i_2 
       (.I0(\custom_alu/MULT [29]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [61]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [29]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[34]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[34]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[19]),
        .I2(CRF_RD2_IBUF[19]),
        .I3(RF_RD2_IBUF[19]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[34]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h5545555555555555)) 
    \Q[34]_i_3 
       (.I0(\Q[30]_i_2__0_n_0 ),
        .I1(EX_CUSTOM_ALU_SEL[28]),
        .I2(EX_CUSTOM_ALU_SEL[26]),
        .I3(EX_CUSTOM_ALU_SEL[27]),
        .I4(\Q[35]_i_7_n_0 ),
        .I5(\Q[34]_i_6_n_0 ),
        .O(\Q[34]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA80AA8080)) 
    \Q[34]_i_3__0 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(\Q[36]_i_3__0_n_0 ),
        .I2(D_MEM_DOUT_IBUF[19]),
        .I3(MEM_D_MEM_ALU_FINAL1),
        .I4(EX_MEM_Q[24]),
        .I5(\Q[36]_i_2__1_n_0 ),
        .O(\Q[34]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'hA8)) 
    \Q[34]_i_4 
       (.I0(\Q[35]_i_11_n_0 ),
        .I1(\Q[35]_i_10_n_0 ),
        .I2(\custom_alu/fp32_mult/exponent_carry__0_n_5 ),
        .O(\Q[34]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \Q[34]_i_5 
       (.I0(EX_CUSTOM_ALU_SEL[30]),
        .I1(EX_CUSTOM_ALU_SEL[29]),
        .I2(EX_CUSTOM_ALU_SEL[31]),
        .O(\Q[34]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h8A800000)) 
    \Q[34]_i_6 
       (.I0(\Q[35]_i_8_n_0 ),
        .I1(ID_EX_Q[126]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(EX_RF_RD1[0]),
        .I4(\Q[35]_i_9_n_0 ),
        .O(\Q[34]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[35]_i_1 
       (.I0(\Q[35]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[20]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[20]),
        .I5(\Q[35]_i_3__0_n_0 ),
        .O(ID_RD2_FORWARDED[20]));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \Q[35]_i_10 
       (.I0(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .I1(\Q[69]_i_14_n_0 ),
        .I2(\Q[69]_i_13_n_0 ),
        .O(\Q[35]_i_10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT5 #(
    .INIT(32'h00000070)) 
    \Q[35]_i_11 
       (.I0(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .I1(\custom_alu/fp32_mult/p_0_in1_in ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\Q[69]_i_14_n_0 ),
        .I4(\Q[69]_i_13_n_0 ),
        .O(\Q[35]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_16 
       (.I0(\custom_alu/int2fp/INT_VAL0 [28]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[154]),
        .I5(EX_RF_RD1[28]),
        .O(\Q[35]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_17 
       (.I0(\custom_alu/int2fp/INT_VAL0 [27]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[153]),
        .I5(EX_RF_RD1[27]),
        .O(\Q[35]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_18 
       (.I0(\custom_alu/int2fp/INT_VAL0 [29]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[155]),
        .I5(EX_RF_RD1[29]),
        .O(\Q[35]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_19 
       (.I0(\custom_alu/int2fp/INT_VAL0 [11]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[137]),
        .I5(EX_RF_RD1[11]),
        .O(\Q[35]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h8AFF8A00)) 
    \Q[35]_i_1__0 
       (.I0(\Q[35]_i_2_n_0 ),
        .I1(\Q[35]_i_3_n_0 ),
        .I2(\Q[35]_i_4_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[30]),
        .O(data0[30]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[35]_i_1__1 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[35]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[30]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[30]));
  LUT6 #(
    .INIT(64'hFFFFFB0B0000FB0B)) 
    \Q[35]_i_2 
       (.I0(\custom_alu/Q [30]),
        .I1(EX_CUSTOM_ALU_SEL[29]),
        .I2(EX_CUSTOM_ALU_SEL[30]),
        .I3(\custom_alu/MULT [62]),
        .I4(EX_CUSTOM_ALU_SEL[31]),
        .I5(\custom_alu/MULT [30]),
        .O(\Q[35]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_20 
       (.I0(\custom_alu/int2fp/INT_VAL0 [12]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[138]),
        .I5(EX_RF_RD1[12]),
        .O(\Q[35]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_21 
       (.I0(\custom_alu/int2fp/INT_VAL0 [10]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[136]),
        .I5(EX_RF_RD1[10]),
        .O(\Q[35]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_22 
       (.I0(\custom_alu/int2fp/INT_VAL0 [9]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[135]),
        .I5(EX_RF_RD1[9]),
        .O(\Q[35]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFE200E2)) 
    \Q[35]_i_23 
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[142]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [16]),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[35]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \Q[35]_i_24 
       (.I0(ALU_DIN1[14]),
        .I1(\custom_alu/int2fp/INT_VAL0 [14]),
        .I2(ALU_DIN1[13]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [13]),
        .O(\Q[35]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEA)) 
    \Q[35]_i_25 
       (.I0(\Q[35]_i_32_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [1]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN1[1]),
        .I4(\Q[29]_i_18__0_n_0 ),
        .I5(\Q[17]_i_15_n_0 ),
        .O(\Q[35]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_26 
       (.I0(\custom_alu/int2fp/INT_VAL0 [7]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[133]),
        .I5(EX_RF_RD1[7]),
        .O(\Q[35]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_27 
       (.I0(\custom_alu/int2fp/INT_VAL0 [8]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[134]),
        .I5(EX_RF_RD1[8]),
        .O(\Q[35]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_28 
       (.I0(\custom_alu/int2fp/INT_VAL0 [5]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[131]),
        .I5(EX_RF_RD1[5]),
        .O(\Q[35]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_29 
       (.I0(\custom_alu/int2fp/INT_VAL0 [6]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[132]),
        .I5(EX_RF_RD1[6]),
        .O(\Q[35]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[35]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[20]),
        .I2(CRF_RD2_IBUF[20]),
        .I3(RF_RD2_IBUF[20]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[35]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7F00FFFF)) 
    \Q[35]_i_3 
       (.I0(\Q[35]_i_7_n_0 ),
        .I1(\Q[35]_i_8_n_0 ),
        .I2(\Q[35]_i_9_n_0 ),
        .I3(\Q[30]_i_5_n_0 ),
        .I4(\Q[34]_i_5_n_0 ),
        .I5(\Q[30]_i_2__0_n_0 ),
        .O(\Q[35]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[35]_i_32 
       (.I0(\custom_alu/int2fp/INT_VAL0 [2]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[128]),
        .I5(EX_RF_RD1[2]),
        .O(\Q[35]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_35 
       (.I0(EX_RF_RD1[12]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[138]),
        .O(\Q[35]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_36 
       (.I0(EX_RF_RD1[11]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[137]),
        .O(\Q[35]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_37 
       (.I0(EX_RF_RD1[10]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[136]),
        .O(\Q[35]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_38 
       (.I0(EX_RF_RD1[9]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[135]),
        .O(\Q[35]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_39 
       (.I0(EX_RF_RD1[16]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[142]),
        .O(\Q[35]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA80AA8080)) 
    \Q[35]_i_3__0 
       (.I0(\Q[46]_i_4_n_0 ),
        .I1(\Q[36]_i_3__0_n_0 ),
        .I2(D_MEM_DOUT_IBUF[20]),
        .I3(MEM_D_MEM_ALU_FINAL1),
        .I4(EX_MEM_Q[25]),
        .I5(\Q[36]_i_2__1_n_0 ),
        .O(\Q[35]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'h1F)) 
    \Q[35]_i_4 
       (.I0(\Q[35]_i_10_n_0 ),
        .I1(\custom_alu/fp32_mult/p_0_in1_in ),
        .I2(\Q[35]_i_11_n_0 ),
        .O(\Q[35]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_40 
       (.I0(EX_RF_RD1[15]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[141]),
        .O(\Q[35]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_41 
       (.I0(EX_RF_RD1[14]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[140]),
        .O(\Q[35]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_42 
       (.I0(EX_RF_RD1[13]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[139]),
        .O(\Q[35]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_43 
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[126]),
        .O(\custom_alu/int2fp/INT_VAL1 [0]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_44 
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[130]),
        .O(\custom_alu/int2fp/INT_VAL1 [4]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_45 
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[129]),
        .O(\custom_alu/int2fp/INT_VAL1 [3]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_46 
       (.I0(EX_RF_RD1[2]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[128]),
        .O(\custom_alu/int2fp/INT_VAL1 [2]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_47 
       (.I0(EX_RF_RD1[1]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[127]),
        .O(\custom_alu/int2fp/INT_VAL1 [1]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_48 
       (.I0(EX_RF_RD1[8]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[134]),
        .O(\Q[35]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_49 
       (.I0(EX_RF_RD1[7]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[133]),
        .O(\custom_alu/int2fp/INT_VAL1 [7]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_50 
       (.I0(EX_RF_RD1[6]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[132]),
        .O(\custom_alu/int2fp/INT_VAL1 [6]));
  LUT3 #(
    .INIT(8'h1D)) 
    \Q[35]_i_51 
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(ID_EX_Q[131]),
        .O(\custom_alu/int2fp/INT_VAL1 [5]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \Q[35]_i_7 
       (.I0(\Q[31]_i_7__0_n_0 ),
        .I1(\Q[35]_i_16_n_0 ),
        .I2(\Q[35]_i_17_n_0 ),
        .I3(\Q[29]_i_7_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .I5(\Q[35]_i_18_n_0 ),
        .O(\Q[35]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \Q[35]_i_8 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[35]_i_20_n_0 ),
        .I2(\Q[35]_i_21_n_0 ),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[35]_i_23_n_0 ),
        .I5(\Q[35]_i_24_n_0 ),
        .O(\Q[35]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \Q[35]_i_9 
       (.I0(\Q[35]_i_25_n_0 ),
        .I1(\Q[35]_i_26_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[35]_i_28_n_0 ),
        .I4(\Q[35]_i_29_n_0 ),
        .O(\Q[35]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[36]_i_1 
       (.I0(\Q[36]_i_2__0_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[21]),
        .I3(data1[21]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[21]));
  LUT6 #(
    .INIT(64'hBBBBBBB8B8B8B8B8)) 
    \Q[36]_i_1__0 
       (.I0(CUSTOM_ALU_OUT[31]),
        .I1(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I2(\D_MEM_ADDR_OBUF[31]_inst_i_2_n_0 ),
        .I3(\D_MEM_ADDR_OBUF[31]_inst_i_3_n_0 ),
        .I4(\D_MEM_ADDR_OBUF[31]_inst_i_4_n_0 ),
        .I5(\D_MEM_ADDR_OBUF[30]_inst_i_7_n_0 ),
        .O(data0[31]));
  LUT6 #(
    .INIT(64'hFFFFEAEEEAEEEAEE)) 
    \Q[36]_i_1__1 
       (.I0(\Q[36]_i_2__1_n_0 ),
        .I1(EX_MEM_Q[36]),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(D_MEM_DOUT_IBUF[31]),
        .I5(\Q[36]_i_3__0_n_0 ),
        .O(data1[31]));
  LUT6 #(
    .INIT(64'hFFFBFBFBAAAAAAAA)) 
    \Q[36]_i_2 
       (.I0(\Q[36]_i_3_n_0 ),
        .I1(\Q[36]_i_4_n_0 ),
        .I2(\Q[30]_i_2__0_n_0 ),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\Q[30]_i_5_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[31]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[36]_i_2__0 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[21]),
        .I2(CRF_RD2_IBUF[21]),
        .I3(RF_RD2_IBUF[21]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[36]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0D00080008000800)) 
    \Q[36]_i_2__1 
       (.I0(MEM_LOAD_SEL[6]),
        .I1(\Q[19]_i_2__2_n_0 ),
        .I2(EX_MEM_Q[37]),
        .I3(EX_MEM_Q[39]),
        .I4(MEM_LOAD_SEL[5]),
        .I5(\Q[20]_i_2__2_n_0 ),
        .O(\Q[36]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[36]_i_3 
       (.I0(\custom_alu/MULT [31]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [63]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [31]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[36]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \Q[36]_i_3__0 
       (.I0(MEM_LOAD_SEL[1]),
        .I1(MEM_LOAD_SEL[2]),
        .I2(MEM_D_MEM_ALU_FINAL1),
        .I3(MEM_LOAD_SEL[6]),
        .I4(MEM_LOAD_SEL[5]),
        .I5(\Q[36]_i_4__0_n_0 ),
        .O(\Q[36]_i_3__0_n_0 ));
  LUT4 #(
    .INIT(16'hEBFF)) 
    \Q[36]_i_4 
       (.I0(\Q[69]_i_14_n_0 ),
        .I1(\custom_alu/fp32_mult/a_Q ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[31] ),
        .I3(EX_CUSTOM_ALU_SEL[28]),
        .O(\Q[36]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \Q[36]_i_4__0 
       (.I0(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I1(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .O(\Q[36]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[37]_i_1 
       (.I0(\Q[37]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[22]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[22]),
        .I5(\Q[37]_i_3_n_0 ),
        .O(ID_RD2_FORWARDED[22]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[37]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[22]),
        .I2(CRF_RD2_IBUF[22]),
        .I3(RF_RD2_IBUF[22]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[37]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \Q[37]_i_3 
       (.I0(DIN2_FORWARD[0]),
        .I1(DIN2_FORWARD[1]),
        .I2(data1[22]),
        .O(\Q[37]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[38]_i_1 
       (.I0(\Q[38]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[23]),
        .I3(data1[23]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[23]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[38]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[23]),
        .I2(CRF_RD2_IBUF[23]),
        .I3(RF_RD2_IBUF[23]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[38]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[39]_i_1 
       (.I0(\Q[39]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[24]),
        .I3(data1[24]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[24]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[39]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[24]),
        .I2(CRF_RD2_IBUF[24]),
        .I3(RF_RD2_IBUF[24]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[39]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[3]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [2]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [3]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [3]));
  LUT4 #(
    .INIT(16'h00A8)) 
    \Q[3]_i_1__0 
       (.I0(\Q[3]_i_2_n_0 ),
        .I1(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[4] ),
        .I2(\Q[30]_i_2__1_n_0 ),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [3]));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[3]_i_1__1 
       (.I0(I_MEM_DOUT_IBUF[10]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[10]));
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT5 #(
    .INIT(32'h007F0080)) 
    \Q[3]_i_1__2 
       (.I0(STALL_COUNTER_Q[2]),
        .I1(STALL_COUNTER_Q[0]),
        .I2(STALL_COUNTER_Q[1]),
        .I3(STALL_COUNTER_D1),
        .I4(STALL_COUNTER_Q[3]),
        .O(STALL_COUNTER_D[3]));
  LUT6 #(
    .INIT(64'hF377FFFFF3773333)) 
    \Q[3]_i_2 
       (.I0(\Q[3]_i_3_n_0 ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [23]),
        .I4(\custom_alu/fp32_add/sel0 [24]),
        .I5(\custom_alu/fp32_add/data23 [3]),
        .O(\Q[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4744477747774777)) 
    \Q[3]_i_3 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [20]),
        .O(\Q[3]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[40]_i_1 
       (.I0(\Q[40]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[25]),
        .I3(data1[25]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[25]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[40]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[25]),
        .I2(CRF_RD2_IBUF[25]),
        .I3(RF_RD2_IBUF[25]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[40]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[41]_i_1 
       (.I0(\Q[41]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[26]),
        .I3(data1[26]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[26]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[41]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[26]),
        .I2(CRF_RD2_IBUF[26]),
        .I3(RF_RD2_IBUF[26]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[41]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[42]_i_1 
       (.I0(\Q[42]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[27]),
        .I3(data1[27]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[27]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[42]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[27]),
        .I2(CRF_RD2_IBUF[27]),
        .I3(RF_RD2_IBUF[27]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[42]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[43]_i_1 
       (.I0(\Q[43]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[28]),
        .I3(data1[28]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[28]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[43]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[28]),
        .I2(CRF_RD2_IBUF[28]),
        .I3(RF_RD2_IBUF[28]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[43]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[44]_i_1 
       (.I0(\Q[44]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[29]),
        .I3(data1[29]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[29]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[44]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[29]),
        .I2(CRF_RD2_IBUF[29]),
        .I3(RF_RD2_IBUF[29]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[44]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[45]_i_1 
       (.I0(\Q[45]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[30]),
        .I3(data1[30]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[30]));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[45]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[30]),
        .I2(CRF_RD2_IBUF[30]),
        .I3(RF_RD2_IBUF[30]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[45]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[46]_i_1 
       (.I0(\Q[46]_i_2_n_0 ),
        .I1(\Q[46]_i_3_n_0 ),
        .I2(data0[31]),
        .I3(data1[31]),
        .I4(\Q[46]_i_4_n_0 ),
        .O(ID_RD2_FORWARDED[31]));
  LUT5 #(
    .INIT(32'hFFFF6FF6)) 
    \Q[46]_i_10 
       (.I0(CUSTOM_RS2),
        .I1(WB_CUSTOM_RD),
        .I2(CRF_RA2_OBUF[3]),
        .I3(CRF_WA_OBUF[3]),
        .I4(\Q[46]_i_17_n_0 ),
        .O(\Q[46]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hEFFE)) 
    \Q[46]_i_11 
       (.I0(\Q[46]_i_14_n_0 ),
        .I1(\Q[77]_i_6_n_0 ),
        .I2(CUSTOM_RS2),
        .I3(MEM_CUSTOM_RD),
        .O(\Q[46]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \Q[46]_i_12 
       (.I0(CRF_RA2_OBUF[2]),
        .I1(EX_MEM_Q[2]),
        .I2(CRF_RA2_OBUF[3]),
        .I3(EX_MEM_Q[3]),
        .I4(EX_MEM_Q[4]),
        .I5(CRF_RA2_OBUF[4]),
        .O(\Q[46]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \Q[46]_i_13 
       (.I0(CRF_RA2_OBUF[2]),
        .I1(CRF_WA_OBUF[2]),
        .I2(CRF_RA2_OBUF[0]),
        .I3(CRF_WA_OBUF[0]),
        .I4(CRF_WA_OBUF[1]),
        .I5(CRF_RA2_OBUF[1]),
        .O(\Q[46]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h6FF6)) 
    \Q[46]_i_14 
       (.I0(EX_MEM_Q[1]),
        .I1(CRF_RA2_OBUF[1]),
        .I2(EX_MEM_Q[0]),
        .I3(CRF_RA2_OBUF[0]),
        .O(\Q[46]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hBEFFFFBE)) 
    \Q[46]_i_15 
       (.I0(\Q[78]_i_17_n_0 ),
        .I1(CRF_RA2_OBUF[2]),
        .I2(ID_EX_Q[2]),
        .I3(ID_EX_Q[0]),
        .I4(CRF_RA2_OBUF[0]),
        .O(\Q[46]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h6FF6)) 
    \Q[46]_i_16 
       (.I0(ID_EX_Q[3]),
        .I1(CRF_RA2_OBUF[3]),
        .I2(ID_EX_Q[1]),
        .I3(CRF_RA2_OBUF[1]),
        .O(\Q[46]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hF6)) 
    \Q[46]_i_17 
       (.I0(CRF_WA_OBUF[4]),
        .I1(CRF_RA2_OBUF[4]),
        .I2(\Q[78]_i_15_n_0 ),
        .O(\Q[46]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[46]_i_2 
       (.I0(DIN2_FORWARD[2]),
        .I1(CRF_WD_OBUF[31]),
        .I2(CRF_RD2_IBUF[31]),
        .I3(RF_RD2_IBUF[31]),
        .I4(CUSTOM_RS2),
        .I5(\Q[46]_i_7_n_0 ),
        .O(\Q[46]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \Q[46]_i_3 
       (.I0(\Q[46]_i_7_n_0 ),
        .I1(DIN2_FORWARD[0]),
        .O(\Q[46]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[46]_i_4 
       (.I0(DIN2_FORWARD[1]),
        .I1(DIN2_FORWARD[0]),
        .O(\Q[46]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00005554)) 
    \Q[46]_i_5 
       (.I0(\Q[46]_i_10_n_0 ),
        .I1(\Q[46]_i_11_n_0 ),
        .I2(DIN2_FORWARD[0]),
        .I3(\Q[46]_i_12_n_0 ),
        .I4(\Q[46]_i_13_n_0 ),
        .O(DIN2_FORWARD[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000008)) 
    \Q[46]_i_6 
       (.I0(\Q[0]_i_3_n_0 ),
        .I1(I_MEM_DOUT_IBUF[13]),
        .I2(I_MEM_DOUT_IBUF[12]),
        .I3(I_MEM_DOUT_IBUF[14]),
        .I4(\Q[161]_i_4_n_0 ),
        .I5(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .O(CUSTOM_RS2));
  LUT6 #(
    .INIT(64'hFFFFFFFF01000001)) 
    \Q[46]_i_7 
       (.I0(\Q[46]_i_12_n_0 ),
        .I1(\Q[46]_i_14_n_0 ),
        .I2(\Q[77]_i_6_n_0 ),
        .I3(CUSTOM_RS2),
        .I4(MEM_CUSTOM_RD),
        .I5(DIN2_FORWARD[0]),
        .O(\Q[46]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h1001000000001001)) 
    \Q[46]_i_8 
       (.I0(\Q[46]_i_15_n_0 ),
        .I1(\Q[46]_i_16_n_0 ),
        .I2(EX_CUSTOM_RD),
        .I3(CUSTOM_RS2),
        .I4(ID_EX_Q[4]),
        .I5(CRF_RA2_OBUF[4]),
        .O(DIN2_FORWARD[0]));
  LUT6 #(
    .INIT(64'h0000000000000009)) 
    \Q[46]_i_9 
       (.I0(MEM_CUSTOM_RD),
        .I1(CUSTOM_RS2),
        .I2(\Q[77]_i_6_n_0 ),
        .I3(\Q[46]_i_14_n_0 ),
        .I4(DIN2_FORWARD[0]),
        .I5(\Q[46]_i_12_n_0 ),
        .O(DIN2_FORWARD[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[47]_i_1 
       (.I0(\Q[47]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[0]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[0]),
        .I5(\Q[47]_i_4_n_0 ),
        .O(\Q[47]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[47]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[0]),
        .I2(CRF_RD1_IBUF[0]),
        .I3(RF_RD1_IBUF[0]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[47]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFABAAAAAAAAAA)) 
    \Q[47]_i_3 
       (.I0(\Q[5]_i_2__0_n_0 ),
        .I1(\custom_alu/fp2int/p_0_in [0]),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(EX_CUSTOM_ALU_SEL[27]),
        .I4(\Q[47]_i_5_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[0]));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[47]_i_4 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[0]),
        .O(\Q[47]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF44F444444444)) 
    \Q[47]_i_5 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [0]),
        .I2(\Q[26]_i_7_n_0 ),
        .I3(\Q[47]_i_6_n_0 ),
        .I4(\Q[47]_i_7_n_0 ),
        .I5(\Q[30]_i_5_n_0 ),
        .O(\Q[47]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A888AAA8AAA8AAA)) 
    \Q[47]_i_6 
       (.I0(\Q[47]_i_8_n_0 ),
        .I1(\Q[9]_i_11_n_0 ),
        .I2(\Q[47]_i_9_n_0 ),
        .I3(\Q[29]_i_10_n_0 ),
        .I4(\Q[28]_i_20_n_0 ),
        .I5(ALU_DIN1[0]),
        .O(\Q[47]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[47]_i_7 
       (.I0(\Q[35]_i_26_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[35]_i_29_n_0 ),
        .I4(\Q[35]_i_28_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[47]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000535FFFFF535F)) 
    \Q[47]_i_8 
       (.I0(\Q[29]_i_18__0_n_0 ),
        .I1(\Q[35]_i_32_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[23]_i_13__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[17]_i_15_n_0 ),
        .O(\Q[47]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[47]_i_9 
       (.I0(\custom_alu/int2fp/INT_VAL0 [1]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[127]),
        .I5(EX_RF_RD1[1]),
        .O(\Q[47]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[48]_i_1 
       (.I0(\Q[48]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[1]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[1]),
        .I5(\Q[48]_i_4_n_0 ),
        .O(\Q[48]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0F77)) 
    \Q[48]_i_10 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(ALU_DIN1[0]),
        .I2(\Q[47]_i_9_n_0 ),
        .I3(\Q[28]_i_20_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[48]_i_12_n_0 ),
        .O(\Q[48]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFF54045404)) 
    \Q[48]_i_11 
       (.I0(\Q[29]_i_18__0_n_0 ),
        .I1(ALU_DIN1[25]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(\custom_alu/int2fp/INT_VAL0 [25]),
        .I4(\Q[17]_i_15_n_0 ),
        .I5(\Q[28]_i_12_n_0 ),
        .O(\Q[48]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hEFEAAFAAEAEAAAAA)) 
    \Q[48]_i_12 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\custom_alu/int2fp/INT_VAL0 [24]),
        .I2(PSUM3__0_carry__0_i_10__2_n_0),
        .I3(ALU_DIN1[24]),
        .I4(\custom_alu/int2fp/INT_VAL0 [2]),
        .I5(ALU_DIN1[2]),
        .O(\Q[48]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[48]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[1]),
        .I2(CRF_RD1_IBUF[1]),
        .I3(RF_RD1_IBUF[1]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[48]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[48]_i_3 
       (.I0(\Q[48]_i_5_n_0 ),
        .I1(\Q[65]_i_5_n_0 ),
        .I2(\custom_alu/fp32_mult/product_mantissa [1]),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\Q[48]_i_6_n_0 ),
        .O(CUSTOM_ALU_OUT[1]));
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[48]_i_4 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[1]),
        .O(\Q[48]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0D0D0D0D000D0D0D)) 
    \Q[48]_i_5 
       (.I0(\Q[14]_i_4__0_n_0 ),
        .I1(INT0_carry_i_13_n_0),
        .I2(\Q[48]_i_7_n_0 ),
        .I3(\Q[48]_i_8_n_0 ),
        .I4(\Q[27]_i_7_n_0 ),
        .I5(\Q[48]_i_9_n_0 ),
        .O(\Q[48]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB8B8888BB8B)) 
    \Q[48]_i_6 
       (.I0(\custom_alu/MULT [1]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(EX_CUSTOM_ALU_SEL[29]),
        .I3(\custom_alu/Q [1]),
        .I4(EX_CUSTOM_ALU_SEL[30]),
        .I5(\custom_alu/MULT [33]),
        .O(\Q[48]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[48]_i_7 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [1]),
        .O(\Q[48]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0EFEFFFFFFFFFFFF)) 
    \Q[48]_i_8 
       (.I0(\Q[48]_i_10_n_0 ),
        .I1(\Q[48]_i_11_n_0 ),
        .I2(\Q[35]_i_17_n_0 ),
        .I3(\Q[35]_i_28_n_0 ),
        .I4(\Q[26]_i_7_n_0 ),
        .I5(\Q[27]_i_13_n_0 ),
        .O(\Q[48]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[48]_i_9 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[35]_i_29_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[48]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[49]_i_1 
       (.I0(\Q[49]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[2]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[2]),
        .I5(\Q[49]_i_4_n_0 ),
        .O(\Q[49]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[49]_i_10 
       (.I0(\Q[35]_i_22_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[35]_i_26_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[49]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[49]_i_11 
       (.I0(\Q_reg[49]_i_17_n_6 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_17_n_7 ),
        .O(\Q[49]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[49]_i_12 
       (.I0(\Q_reg[49]_i_18_n_7 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_17_n_4 ),
        .O(\Q[49]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[49]_i_13 
       (.I0(\Q_reg[49]_i_17_n_4 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_17_n_5 ),
        .O(\Q[49]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[49]_i_14 
       (.I0(\Q_reg[49]_i_17_n_5 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_17_n_6 ),
        .O(\Q[49]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h59AA0CF359AAFF00)) 
    \Q[49]_i_15 
       (.I0(\Q_reg[49]_i_17_n_6 ),
        .I1(\Q[49]_i_19_n_0 ),
        .I2(\Q[49]_i_20_n_0 ),
        .I3(\Q_reg[49]_i_17_n_7 ),
        .I4(\custom_alu/fp32_mult/normalised ),
        .I5(\Q_reg[49]_i_21_n_4 ),
        .O(\Q[49]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FF07)) 
    \Q[49]_i_16 
       (.I0(\Q[31]_i_14__0_n_0 ),
        .I1(ALU_DIN1[0]),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[49]_i_22_n_0 ),
        .I4(\Q[29]_i_7_n_0 ),
        .I5(\Q[49]_i_23_n_0 ),
        .O(\Q[49]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \Q[49]_i_19 
       (.I0(\custom_alu/fp32_mult/p_1_in [3]),
        .I1(\custom_alu/fp32_mult/p_1_in [9]),
        .I2(\Q_reg[49]_i_32_n_6 ),
        .I3(\Q_reg[49]_i_21_n_7 ),
        .I4(\Q[49]_i_33_n_0 ),
        .O(\Q[49]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[49]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[2]),
        .I2(CRF_RD1_IBUF[2]),
        .I3(RF_RD1_IBUF[2]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[49]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \Q[49]_i_20 
       (.I0(\Q[49]_i_34_n_0 ),
        .I1(\Q_reg[49]_i_21_n_5 ),
        .I2(\Q_reg[49]_i_35_n_5 ),
        .I3(\custom_alu/fp32_mult/p_1_in [10]),
        .I4(\custom_alu/fp32_mult/p_1_in [5]),
        .I5(\Q[49]_i_36_n_0 ),
        .O(\Q[49]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h000004F4FFFF04F4)) 
    \Q[49]_i_22 
       (.I0(\Q[47]_i_9_n_0 ),
        .I1(\Q[31]_i_13__0_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[35]_i_32_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[29]_i_18__0_n_0 ),
        .O(\Q[49]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h5555555533300030)) 
    \Q[49]_i_23 
       (.I0(\Q[35]_i_28_n_0 ),
        .I1(\Q[17]_i_15_n_0 ),
        .I2(ALU_DIN1[25]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [25]),
        .I5(\Q[28]_i_12_n_0 ),
        .O(\Q[49]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[49]_i_3 
       (.I0(\Q[49]_i_5_n_0 ),
        .I1(\Q[65]_i_5_n_0 ),
        .I2(\custom_alu/fp32_mult/product_mantissa [2]),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\Q[49]_i_7_n_0 ),
        .O(CUSTOM_ALU_OUT[2]));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \Q[49]_i_33 
       (.I0(\Q_reg[49]_i_21_n_4 ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\Q_reg[49]_i_32_n_4 ),
        .I3(\Q_reg[49]_i_32_n_7 ),
        .O(\Q[49]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \Q[49]_i_34 
       (.I0(\Q_reg[49]_i_21_n_6 ),
        .I1(\Q_reg[49]_i_35_n_4 ),
        .I2(\Q_reg[49]_i_35_n_7 ),
        .I3(\custom_alu/fp32_mult/p_1_in [1]),
        .O(\Q[49]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \Q[49]_i_36 
       (.I0(\custom_alu/fp32_mult/p_1_in [7]),
        .I1(\Q_reg[49]_i_32_n_5 ),
        .I2(\custom_alu/fp32_mult/p_1_in [2]),
        .I3(\Q_reg[49]_i_35_n_6 ),
        .I4(\Q[49]_i_48_n_0 ),
        .O(\Q[49]_i_36_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[49]_i_4 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[2]),
        .O(\Q[49]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \Q[49]_i_48 
       (.I0(\custom_alu/fp32_mult/p_1_in [8]),
        .I1(\custom_alu/fp32_mult/p_1_in [4]),
        .I2(\custom_alu/fp32_mult/p_1_in [6]),
        .I3(\custom_alu/fp32_mult/p_1_in [0]),
        .O(\Q[49]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0D0D0D0D000D0D0D)) 
    \Q[49]_i_5 
       (.I0(\Q[14]_i_4__0_n_0 ),
        .I1(INT0_carry_i_12_n_0),
        .I2(\Q[49]_i_8_n_0 ),
        .I3(\Q[49]_i_9_n_0 ),
        .I4(\Q[27]_i_7_n_0 ),
        .I5(\Q[49]_i_10_n_0 ),
        .O(\Q[49]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB8B8888BB8B)) 
    \Q[49]_i_7 
       (.I0(\custom_alu/MULT [2]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(EX_CUSTOM_ALU_SEL[29]),
        .I3(\custom_alu/Q [2]),
        .I4(EX_CUSTOM_ALU_SEL[30]),
        .I5(\custom_alu/MULT [34]),
        .O(\Q[49]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[49]_i_8 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [2]),
        .O(\Q[49]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h2EFFFFFF)) 
    \Q[49]_i_9 
       (.I0(\Q[49]_i_16_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[35]_i_29_n_0 ),
        .I3(\Q[26]_i_7_n_0 ),
        .I4(\Q[27]_i_13_n_0 ),
        .O(\Q[49]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT4 #(
    .INIT(16'h0B08)) 
    \Q[4]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [4]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\Q[30]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/significand_add0 [3]),
        .O(\custom_alu/fp32_add/p_1_out [4]));
  LUT3 #(
    .INIT(8'h5C)) 
    \Q[4]_i_11 
       (.I0(\Q[8]_i_13_n_0 ),
        .I1(\Q[4]_i_20_n_0 ),
        .I2(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[4]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[4]_i_12 
       (.I0(\Q[12]_i_19_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[8]_i_18_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[4]_i_15_n_0 ),
        .O(\Q[4]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \Q[4]_i_13 
       (.I0(\Q[4]_i_20_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\Q[8]_i_17_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I4(\Q[4]_i_21_n_0 ),
        .O(\Q[4]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \Q[4]_i_14 
       (.I0(\Q[8]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[4]_i_22_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I4(\Q[4]_i_23_n_0 ),
        .O(\Q[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \Q[4]_i_15 
       (.I0(\Q[8]_i_16_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[4]_i_24_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I4(\Q[4]_i_25_n_0 ),
        .O(\Q[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \Q[4]_i_16 
       (.I0(ALU_DIN2[3]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[129]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[3]),
        .O(\Q[4]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \Q[4]_i_17 
       (.I0(ALU_DIN2[2]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[128]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[2]),
        .O(\Q[4]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \Q[4]_i_18 
       (.I0(ALU_DIN2[1]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[127]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[1]),
        .O(\Q[4]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \Q[4]_i_19 
       (.I0(\Q[23]_i_13_n_0 ),
        .I1(\Q[4]_i_15_n_0 ),
        .I2(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I3(\Q[4]_i_14_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [0]),
        .O(\Q[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[4]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[5] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/data23 [4]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\Q[4]_i_3__0_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [4]));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[4]_i_1__1 
       (.I0(I_MEM_DOUT_IBUF[11]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[11]));
  LUT6 #(
    .INIT(64'h00007FFF00008000)) 
    \Q[4]_i_1__2 
       (.I0(STALL_COUNTER_Q[3]),
        .I1(STALL_COUNTER_Q[1]),
        .I2(STALL_COUNTER_Q[0]),
        .I3(STALL_COUNTER_Q[2]),
        .I4(STALL_COUNTER_D1),
        .I5(STALL_COUNTER_Q[4]),
        .O(STALL_COUNTER_D[4]));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[4]_i_2 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[4]),
        .I2(STALL_EN),
        .I3(IF_PC2[4]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[4] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[4]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h47444777)) 
    \Q[4]_i_20 
       (.I0(\Q[8]_i_15_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[12]_i_20_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I4(\Q[4]_i_26_n_0 ),
        .O(\Q[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[4]_i_21 
       (.I0(ALU_DIN2[9]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[9]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[4]_i_27_n_0 ),
        .O(\Q[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[4]_i_22 
       (.I0(EX_RF_RD2[8]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[87]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[8]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \Q[4]_i_23 
       (.I0(ALU_DIN1[16]),
        .I1(ALU_DIN2[16]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I3(ALU_DIN1[0]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[0]),
        .O(\Q[4]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[4]_i_24 
       (.I0(EX_RF_RD2[10]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[89]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[10]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(\Q[4]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \Q[4]_i_25 
       (.I0(ALU_DIN1[18]),
        .I1(ALU_DIN2[18]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I3(ALU_DIN1[2]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[2]),
        .O(\Q[4]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \Q[4]_i_26 
       (.I0(ALU_DIN1[19]),
        .I1(ALU_DIN2[19]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I3(ALU_DIN1[3]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[3]),
        .O(\Q[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \Q[4]_i_27 
       (.I0(ALU_DIN1[17]),
        .I1(ALU_DIN2[17]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I3(ALU_DIN1[1]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[1]),
        .O(\Q[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000D1)) 
    \Q[4]_i_3 
       (.I0(\Q[4]_i_11_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[8]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [6]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [7]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \Q[4]_i_3__0 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\Q[4]_i_9_n_0 ),
        .O(\Q[4]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[4]_i_3__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[3]),
        .I2(STALL_EN),
        .I3(IF_PC2[3]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[3] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[4]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000074)) 
    \Q[4]_i_4 
       (.I0(\Q[4]_i_11_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[4]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [6]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [7]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [2]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[4]_i_4__0 
       (.I0(\custom_alu/fp32_add/sel0 [0]),
        .O(\Q[4]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h001BFF1BFFFFFFFF)) 
    \Q[4]_i_4__1 
       (.I0(EX_BR_TAKEN),
        .I1(\FF_IF_ID_PCADD/Q_reg_n_0_[2] ),
        .I2(IF_PC2[2]),
        .I3(STALL_EN),
        .I4(ID_PC[2]),
        .I5(RSTn_IBUF),
        .O(\Q[4]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000D1)) 
    \Q[4]_i_5 
       (.I0(\Q[4]_i_13_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[4]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [6]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [5]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [7]),
        .O(\custom_alu/fp32_add/significand_b_add_sub [1]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[4]_i_5__0 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .O(\Q[4]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[4]_i_5__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[1]),
        .I2(STALL_EN),
        .I3(IF_PC2[1]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[1] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[4]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000077744474)) 
    \Q[4]_i_6 
       (.I0(\Q[4]_i_13_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[4]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[4]_i_15_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [0]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[4]_i_6__0 
       (.I0(\custom_alu/fp32_add/sel0 [3]),
        .O(\Q[4]_i_6__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[4]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .O(\Q[4]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[4]_i_8 
       (.I0(\custom_alu/fp32_add/sel0 [1]),
        .O(\Q[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[4]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [21]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [20]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [19]),
        .O(\Q[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[50]_i_1 
       (.I0(\Q[50]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[3]),
        .I4(data1[3]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[50]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[50]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[3]),
        .I3(CRF_RD1_IBUF[3]),
        .I4(CRF_WD_OBUF[3]),
        .O(\Q[50]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[51]_i_1 
       (.I0(\Q[51]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[4]),
        .I4(data1[4]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[51]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[51]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[4]),
        .I3(CRF_RD1_IBUF[4]),
        .I4(CRF_WD_OBUF[4]),
        .O(\Q[51]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[52]_i_1 
       (.I0(\Q[52]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[5]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[5]),
        .I5(\Q[52]_i_4_n_0 ),
        .O(\Q[52]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[52]_i_10 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_19_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[35]_i_21_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[52]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8888888B888)) 
    \Q[52]_i_11 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[28]_i_12_n_0 ),
        .I2(\Q[35]_i_26_n_0 ),
        .I3(ALU_DIN1[25]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [25]),
        .O(\Q[52]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF4444444F444)) 
    \Q[52]_i_12 
       (.I0(\Q[21]_i_10__0_n_0 ),
        .I1(\Q[47]_i_9_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[35]_i_32_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[29]_i_18__0_n_0 ),
        .O(\Q[52]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000004F4FFFF04F4)) 
    \Q[52]_i_13 
       (.I0(\Q[17]_i_15_n_0 ),
        .I1(\Q[31]_i_13__0_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[35]_i_28_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[35]_i_29_n_0 ),
        .O(\Q[52]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[52]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[5]),
        .I2(CRF_RD1_IBUF[5]),
        .I3(RF_RD1_IBUF[5]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[52]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBBBFBBBBAAAAAAAA)) 
    \Q[52]_i_3 
       (.I0(\Q[10]_i_2__0_n_0 ),
        .I1(\Q[10]_i_3_n_0 ),
        .I2(\Q[52]_i_5_n_0 ),
        .I3(\Q[52]_i_6_n_0 ),
        .I4(\Q[52]_i_7_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[5]));
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[52]_i_4 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(data1[5]),
        .O(\Q[52]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000115155555555)) 
    \Q[52]_i_5 
       (.I0(EX_CUSTOM_ALU_SEL[27]),
        .I1(\Q[26]_i_7_n_0 ),
        .I2(\Q[52]_i_8_n_0 ),
        .I3(\Q[52]_i_9_n_0 ),
        .I4(\Q[52]_i_10_n_0 ),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[52]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[52]_i_6 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__0_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [5]),
        .O(\Q[52]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEFEAFFFF)) 
    \Q[52]_i_7 
       (.I0(INT0_carry__0_i_9_n_0),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__1_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[52]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBAAAB)) 
    \Q[52]_i_8 
       (.I0(\Q[35]_i_17_n_0 ),
        .I1(\Q[52]_i_11_n_0 ),
        .I2(\Q[52]_i_12_n_0 ),
        .I3(\Q[67]_i_12_n_0 ),
        .I4(\Q[52]_i_13_n_0 ),
        .I5(\Q[29]_i_7_n_0 ),
        .O(\Q[52]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFF404040)) 
    \Q[52]_i_9 
       (.I0(\Q[13]_i_11_n_0 ),
        .I1(\Q[28]_i_11_n_0 ),
        .I2(ALU_DIN1[0]),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .O(\Q[52]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[53]_i_1 
       (.I0(\Q[53]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[6]),
        .I4(data1[6]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[53]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[53]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[6]),
        .I3(CRF_RD1_IBUF[6]),
        .I4(CRF_WD_OBUF[6]),
        .O(\Q[53]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[54]_i_1 
       (.I0(\Q[54]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[7]),
        .I4(data1[7]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[54]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[54]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[7]),
        .I3(CRF_RD1_IBUF[7]),
        .I4(CRF_WD_OBUF[7]),
        .O(\Q[54]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[55]_i_1 
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[23]),
        .O(\custom_alu/fp32_add/p_0_in [0]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[55]_i_1__0 
       (.I0(\Q[55]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[8]),
        .I4(data1[8]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[55]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[55]_i_1__1 
       (.I0(ID_EX_Q[149]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[23]),
        .O(ALU_DIN1[23]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[55]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[8]),
        .I3(CRF_RD1_IBUF[8]),
        .I4(CRF_WD_OBUF[8]),
        .O(\Q[55]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[56]_i_1 
       (.I0(ID_EX_Q[103]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[24]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[24]),
        .O(\custom_alu/fp32_add/p_0_in [1]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[56]_i_1__0 
       (.I0(\Q[56]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[9]),
        .I4(data1[9]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[56]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[56]_i_1__1 
       (.I0(ID_EX_Q[150]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[24]),
        .O(ALU_DIN1[24]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[56]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[9]),
        .I3(CRF_RD1_IBUF[9]),
        .I4(CRF_WD_OBUF[9]),
        .O(\Q[56]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[57]_i_1 
       (.I0(ID_EX_Q[104]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[25]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[25]),
        .O(\custom_alu/fp32_add/p_0_in [2]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[57]_i_1__0 
       (.I0(\Q[57]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[10]),
        .I4(data1[10]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[57]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[57]_i_1__1 
       (.I0(ID_EX_Q[151]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[25]),
        .O(ALU_DIN1[25]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[57]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[10]),
        .I3(CRF_RD1_IBUF[10]),
        .I4(CRF_WD_OBUF[10]),
        .O(\Q[57]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[58]_i_1 
       (.I0(ID_EX_Q[105]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[26]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[26]),
        .O(\custom_alu/fp32_add/p_0_in [3]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[58]_i_1__0 
       (.I0(\Q[58]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[11]),
        .I4(data1[11]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[58]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[58]_i_1__1 
       (.I0(ID_EX_Q[152]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[26]),
        .O(ALU_DIN1[26]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[58]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[11]),
        .I3(CRF_RD1_IBUF[11]),
        .I4(CRF_WD_OBUF[11]),
        .O(\Q[58]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[59]_i_1 
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[27]),
        .O(\custom_alu/fp32_add/p_0_in [4]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[59]_i_1__0 
       (.I0(\Q[59]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[12]),
        .I4(data1[12]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[59]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[59]_i_1__1 
       (.I0(ID_EX_Q[153]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[27]),
        .O(ALU_DIN1[27]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[59]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[12]),
        .I3(CRF_RD1_IBUF[12]),
        .I4(CRF_WD_OBUF[12]),
        .O(\Q[59]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[5]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [5]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [4]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [5]));
  LUT5 #(
    .INIT(32'h00000777)) 
    \Q[5]_i_10 
       (.I0(\Q[28]_i_7_n_0 ),
        .I1(\Q[35]_i_28_n_0 ),
        .I2(\Q[35]_i_29_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .O(\Q[5]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[5]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[6] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\Q[5]_i_2_n_0 ),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [5]));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \Q[5]_i_1__1 
       (.I0(\Q[5]_i_2__0_n_0 ),
        .I1(\Q[5]_i_3_n_0 ),
        .I2(\Q[34]_i_5_n_0 ),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(D_MEM_ADDR_OBUF[0]),
        .O(data0[0]));
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \Q[5]_i_1__2 
       (.I0(\Q[5]_i_2__1_n_0 ),
        .I1(\Q[11]_i_3__0_n_0 ),
        .I2(\Q[5]_i_3__1_n_0 ),
        .I3(\Q[11]_i_5__1_n_0 ),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(EX_MEM_Q[5]),
        .O(data1[0]));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'h12)) 
    \Q[5]_i_1__3 
       (.I0(\Q[5]_i_2__2_n_0 ),
        .I1(STALL_COUNTER_D1),
        .I2(STALL_COUNTER_Q[5]),
        .O(STALL_COUNTER_D[5]));
  LUT5 #(
    .INIT(32'h8B8BFF00)) 
    \Q[5]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\Q[5]_i_3__0_n_0 ),
        .I3(\custom_alu/fp32_add/data23 [5]),
        .I4(\custom_alu/fp32_add/sel0 [24]),
        .O(\Q[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[5]_i_2__0 
       (.I0(\custom_alu/MULT [0]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [32]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [0]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[5]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[5]_i_2__1 
       (.I0(D_MEM_DOUT_IBUF[8]),
        .I1(D_MEM_DOUT_IBUF[0]),
        .I2(D_MEM_DOUT_IBUF[24]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[16]),
        .O(\Q[5]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \Q[5]_i_2__2 
       (.I0(STALL_COUNTER_Q[4]),
        .I1(STALL_COUNTER_Q[2]),
        .I2(STALL_COUNTER_Q[0]),
        .I3(STALL_COUNTER_Q[1]),
        .I4(STALL_COUNTER_Q[3]),
        .O(\Q[5]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h00EF00EF000000EF)) 
    \Q[5]_i_3 
       (.I0(\custom_alu/fp2int/p_0_in [0]),
        .I1(EX_CUSTOM_ALU_SEL[28]),
        .I2(EX_CUSTOM_ALU_SEL[27]),
        .I3(\Q[5]_i_5_n_0 ),
        .I4(\custom_alu/fp32_mult/product_mantissa [0]),
        .I5(\Q[65]_i_5_n_0 ),
        .O(\Q[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0047FF47)) 
    \Q[5]_i_3__0 
       (.I0(\custom_alu/fp32_add/sel0 [3]),
        .I1(\custom_alu/fp32_add/sel0 [21]),
        .I2(\Q[5]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [4]),
        .O(\Q[5]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[5]_i_3__1 
       (.I0(D_MEM_DOUT_IBUF[0]),
        .I1(D_MEM_DOUT_IBUF[16]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[24]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[8]),
        .O(\Q[5]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[5]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [20]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [19]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [18]),
        .O(\Q[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000A8080202AA0A)) 
    \Q[5]_i_5 
       (.I0(\Q[30]_i_5_n_0 ),
        .I1(\Q[26]_i_15__0_n_0 ),
        .I2(\Q[28]_i_6_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[5]_i_10_n_0 ),
        .I5(\Q[47]_i_6_n_0 ),
        .O(\Q[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[60]_i_1 
       (.I0(ID_EX_Q[107]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[28]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[28]),
        .O(\custom_alu/fp32_add/p_0_in [5]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[60]_i_1__0 
       (.I0(\Q[60]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[13]),
        .I4(data1[13]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[60]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[60]_i_1__1 
       (.I0(ID_EX_Q[154]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[28]),
        .O(ALU_DIN1[28]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[60]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[13]),
        .I3(CRF_RD1_IBUF[13]),
        .I4(CRF_WD_OBUF[13]),
        .O(\Q[60]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[61]_i_1 
       (.I0(ID_EX_Q[108]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(EX_RF_RD2[29]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[29]),
        .O(\custom_alu/fp32_add/p_0_in [6]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[61]_i_1__0 
       (.I0(\Q[61]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[14]),
        .I4(data1[14]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[61]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[61]_i_1__1 
       (.I0(ID_EX_Q[155]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[29]),
        .O(ALU_DIN1[29]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[61]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[14]),
        .I3(CRF_RD1_IBUF[14]),
        .I4(CRF_WD_OBUF[14]),
        .O(\Q[61]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[62]_i_1 
       (.I0(ID_EX_Q[109]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I2(EX_RF_RD2[30]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[30]),
        .O(\custom_alu/fp32_add/p_0_in [7]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[62]_i_1__0 
       (.I0(\Q[62]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[15]),
        .I4(data1[15]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[62]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[62]_i_1__1 
       (.I0(ID_EX_Q[156]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[30]),
        .O(ALU_DIN1[30]));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[62]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[15]),
        .I3(CRF_RD1_IBUF[15]),
        .I4(CRF_WD_OBUF[15]),
        .O(\Q[62]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[63]_i_1 
       (.I0(\Q[63]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[16]),
        .I4(data1[16]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[63]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[63]_i_1__0 
       (.I0(RSTn_IBUF),
        .O(RST0));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[63]_i_1__1 
       (.I0(ID_EX_Q[157]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I2(EX_RF_RD1[31]),
        .O(\Q[63]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[63]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[16]),
        .I3(CRF_RD1_IBUF[16]),
        .I4(CRF_WD_OBUF[16]),
        .O(\Q[63]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[64]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [0]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [64]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[64]_i_1__0 
       (.I0(\Q[64]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[17]),
        .I4(data1[17]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[64]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[64]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[17]),
        .I3(CRF_RD1_IBUF[17]),
        .I4(CRF_WD_OBUF[17]),
        .O(\Q[64]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[65]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [1]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [65]));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[65]_i_10 
       (.I0(exponent_carry_i_10_n_4),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_10_n_5),
        .O(\Q[65]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[65]_i_11 
       (.I0(exponent_carry_i_10_n_5),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_10_n_6),
        .O(\Q[65]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[65]_i_12 
       (.I0(exponent_carry_i_10_n_6),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_10_n_7),
        .O(\Q[65]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011115155)) 
    \Q[65]_i_13 
       (.I0(\Q[27]_i_13_n_0 ),
        .I1(\Q[69]_i_20_n_0 ),
        .I2(\Q[17]_i_15_n_0 ),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[65]_i_17_n_0 ),
        .I5(\Q[23]_i_14__0_n_0 ),
        .O(\Q[65]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8888888A8A8A888A)) 
    \Q[65]_i_14 
       (.I0(\Q[22]_i_7__0_n_0 ),
        .I1(\Q[65]_i_18_n_0 ),
        .I2(\Q[66]_i_13_n_0 ),
        .I3(\Q[65]_i_19_n_0 ),
        .I4(\Q[35]_i_20_n_0 ),
        .I5(\Q[35]_i_26_n_0 ),
        .O(\Q[65]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFA2)) 
    \Q[65]_i_15 
       (.I0(\Q[65]_i_20_n_0 ),
        .I1(\Q[65]_i_21_n_0 ),
        .I2(\Q[67]_i_12_n_0 ),
        .I3(\Q[29]_i_7_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[65]_i_22_n_0 ),
        .O(\Q[65]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAEEEAE)) 
    \Q[65]_i_16 
       (.I0(INT0_carry_i_6_n_0),
        .I1(INT0_carry__3_i_8_n_0),
        .I2(EX_RF_RD1[23]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I4(ID_EX_Q[149]),
        .I5(INT0_carry__3_i_7_n_0),
        .O(\custom_alu/fp2int/p_0_in [18]));
  LUT6 #(
    .INIT(64'h0000000000FFF4F4)) 
    \Q[65]_i_17 
       (.I0(\Q[35]_i_32_n_0 ),
        .I1(\Q[35]_i_26_n_0 ),
        .I2(\Q[65]_i_23_n_0 ),
        .I3(\Q[29]_i_18__0_n_0 ),
        .I4(\Q[35]_i_27_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[65]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h5555303F55553030)) 
    \Q[65]_i_18 
       (.I0(\Q[35]_i_21_n_0 ),
        .I1(\Q[35]_i_22_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[65]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8888888B888)) 
    \Q[65]_i_19 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_19_n_0 ),
        .I2(\Q[35]_i_28_n_0 ),
        .I3(ALU_DIN1[10]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\custom_alu/int2fp/INT_VAL0 [10]),
        .O(\Q[65]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[65]_i_1__0 
       (.I0(\Q[65]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[18]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[18]),
        .I5(\Q[65]_i_4_n_0 ),
        .O(\Q[65]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[65]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[18]),
        .I2(CRF_RD1_IBUF[18]),
        .I3(RF_RD1_IBUF[18]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[65]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[65]_i_20 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[31]_i_10__0_n_0 ),
        .O(\Q[65]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hF808F808FFFFF808)) 
    \Q[65]_i_21 
       (.I0(\Q[17]_i_14_n_0 ),
        .I1(\Q[31]_i_11__0_n_0 ),
        .I2(\Q[31]_i_14__0_n_0 ),
        .I3(\Q[17]_i_10__0_n_0 ),
        .I4(\Q[17]_i_11__0_n_0 ),
        .I5(\Q[21]_i_10__0_n_0 ),
        .O(\Q[65]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[65]_i_22 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[31]_i_11__0_n_0 ),
        .I5(\Q[23]_i_13__0_n_0 ),
        .O(\Q[65]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h000007F7)) 
    \Q[65]_i_23 
       (.I0(ALU_DIN1[0]),
        .I1(\Q[35]_i_28_n_0 ),
        .I2(\Q[35]_i_29_n_0 ),
        .I3(\Q[47]_i_9_n_0 ),
        .I4(\Q[35]_i_26_n_0 ),
        .O(\Q[65]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFBAAAAAAAAA)) 
    \Q[65]_i_3 
       (.I0(\Q[23]_i_2_n_0 ),
        .I1(\Q[65]_i_5_n_0 ),
        .I2(\custom_alu/fp32_mult/product_mantissa [18]),
        .I3(\Q[65]_i_7_n_0 ),
        .I4(\Q[65]_i_8_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[18]));
  LUT6 #(
    .INIT(64'hAAAAAAAA80AA8080)) 
    \Q[65]_i_4 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(\Q[36]_i_3__0_n_0 ),
        .I2(D_MEM_DOUT_IBUF[18]),
        .I3(MEM_D_MEM_ALU_FINAL1),
        .I4(EX_MEM_Q[23]),
        .I5(\Q[36]_i_2__1_n_0 ),
        .O(\Q[65]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \Q[65]_i_5 
       (.I0(\Q[69]_i_13_n_0 ),
        .I1(\Q[69]_i_14_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .O(\Q[65]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \Q[65]_i_7 
       (.I0(\Q[30]_i_5_n_0 ),
        .I1(\Q[23]_i_6__0_n_0 ),
        .I2(\Q[65]_i_13_n_0 ),
        .I3(\Q[65]_i_14_n_0 ),
        .I4(\Q[65]_i_15_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[65]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h40004050)) 
    \Q[65]_i_8 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(\custom_alu/fp2int/INT0 [18]),
        .I2(EX_CUSTOM_ALU_SEL[27]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/fp2int/p_0_in [18]),
        .O(\Q[65]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[65]_i_9 
       (.I0(exponent_carry_i_9_n_7),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(exponent_carry_i_10_n_4),
        .O(\Q[65]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[66]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [2]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [66]));
  LUT6 #(
    .INIT(64'h5555003F55550000)) 
    \Q[66]_i_10 
       (.I0(\Q[28]_i_20_n_0 ),
        .I1(\Q[28]_i_21_n_0 ),
        .I2(\Q[31]_i_14__0_n_0 ),
        .I3(\Q[66]_i_17_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[66]_i_18_n_0 ),
        .O(\Q[66]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h5555303F55553030)) 
    \Q[66]_i_11 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[35]_i_21_n_0 ),
        .I2(\Q[17]_i_11__0_n_0 ),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[28]_i_18_n_0 ),
        .O(\Q[66]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8888888B888)) 
    \Q[66]_i_12 
       (.I0(\Q[35]_i_26_n_0 ),
        .I1(\Q[35]_i_19_n_0 ),
        .I2(\Q[35]_i_29_n_0 ),
        .I3(ALU_DIN1[10]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(\custom_alu/int2fp/INT_VAL0 [10]),
        .O(\Q[66]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFEFEFF)) 
    \Q[66]_i_13 
       (.I0(\Q[17]_i_11__0_n_0 ),
        .I1(\Q[28]_i_18_n_0 ),
        .I2(\Q[17]_i_14_n_0 ),
        .I3(\Q[35]_i_21_n_0 ),
        .I4(\Q[35]_i_19_n_0 ),
        .I5(\Q[35]_i_20_n_0 ),
        .O(\Q[66]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[66]_i_14 
       (.I0(\Q[35]_i_32_n_0 ),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[47]_i_9_n_0 ),
        .I3(\Q[35]_i_28_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .I5(ALU_DIN1[0]),
        .O(\Q[66]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFC000C0)) 
    \Q[66]_i_15 
       (.I0(\Q[35]_i_28_n_0 ),
        .I1(\Q[35]_i_26_n_0 ),
        .I2(\Q[29]_i_18__0_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[66]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000F44FFFF0F44)) 
    \Q[66]_i_16 
       (.I0(\Q[35]_i_20_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[28]_i_18_n_0 ),
        .I3(\Q[69]_i_16_n_0 ),
        .I4(\Q[28]_i_11_n_0 ),
        .I5(\Q[17]_i_11__0_n_0 ),
        .O(\Q[66]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \Q[66]_i_17 
       (.I0(EX_RF_RD1[22]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[148]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(\custom_alu/int2fp/INT_VAL0 [22]),
        .I5(\Q[28]_i_12_n_0 ),
        .O(\Q[66]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEFAAAAAAAA)) 
    \Q[66]_i_18 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(\Q[67]_i_12_n_0 ),
        .I2(\Q[66]_i_19_n_0 ),
        .I3(\Q[21]_i_10__0_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[66]_i_20_n_0 ),
        .O(\Q[66]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB800B800B800)) 
    \Q[66]_i_19 
       (.I0(\custom_alu/int2fp/INT_VAL0 [17]),
        .I1(PSUM3__0_carry__0_i_10__2_n_0),
        .I2(ALU_DIN1[17]),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[31]_i_11__0_n_0 ),
        .I5(\Q[17]_i_10__0_n_0 ),
        .O(\Q[66]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[66]_i_1__0 
       (.I0(\Q[66]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[19]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[19]),
        .I5(\Q[66]_i_4_n_0 ),
        .O(\Q[66]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[66]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[19]),
        .I2(CRF_RD1_IBUF[19]),
        .I3(RF_RD1_IBUF[19]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[66]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[66]_i_20 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(\Q[28]_i_11_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[31]_i_10__0_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[31]_i_11__0_n_0 ),
        .O(\Q[66]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBBABA)) 
    \Q[66]_i_3 
       (.I0(\Q[24]_i_2_n_0 ),
        .I1(\Q[24]_i_3__1_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\Q[66]_i_5_n_0 ),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\Q[66]_i_6_n_0 ),
        .O(CUSTOM_ALU_OUT[19]));
  LUT6 #(
    .INIT(64'hAAAAAAAA80AA8080)) 
    \Q[66]_i_4 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(\Q[36]_i_3__0_n_0 ),
        .I2(D_MEM_DOUT_IBUF[19]),
        .I3(MEM_D_MEM_ALU_FINAL1),
        .I4(EX_MEM_Q[24]),
        .I5(\Q[36]_i_2__1_n_0 ),
        .O(\Q[66]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h02A20000FEAE0000)) 
    \Q[66]_i_5 
       (.I0(\custom_alu/fp2int/p_0_in [19]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [19]),
        .O(\Q[66]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \Q[66]_i_6 
       (.I0(EX_CUSTOM_ALU_SEL[26]),
        .I1(\Q[66]_i_7_n_0 ),
        .I2(\Q[66]_i_8_n_0 ),
        .I3(\Q[66]_i_9_n_0 ),
        .I4(\Q[66]_i_10_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[66]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[66]_i_7 
       (.I0(\Q[28]_i_12_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[23]_i_13__0_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[66]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h55555404FFFFFFFF)) 
    \Q[66]_i_8 
       (.I0(\Q[66]_i_11_n_0 ),
        .I1(\Q[66]_i_12_n_0 ),
        .I2(\Q[35]_i_20_n_0 ),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[66]_i_13_n_0 ),
        .I5(\Q[22]_i_7__0_n_0 ),
        .O(\Q[66]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4700)) 
    \Q[66]_i_9 
       (.I0(\Q[66]_i_14_n_0 ),
        .I1(\Q[69]_i_22_n_0 ),
        .I2(\Q[66]_i_15_n_0 ),
        .I3(\Q[69]_i_20_n_0 ),
        .I4(\Q[66]_i_16_n_0 ),
        .I5(\Q[27]_i_13_n_0 ),
        .O(\Q[66]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[67]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [3]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [67]));
  LUT5 #(
    .INIT(32'hAA8A888A)) 
    \Q[67]_i_10 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[4]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[4]_i_11_n_0 ),
        .O(\Q[67]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000535FFFFF535F)) 
    \Q[67]_i_10__0 
       (.I0(\Q[28]_i_20_n_0 ),
        .I1(\Q[31]_i_13__0_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[23]_i_13__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[29]_i_10_n_0 ),
        .O(\Q[67]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'h8AAA8A88)) 
    \Q[67]_i_11 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[4]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[4]_i_13_n_0 ),
        .O(\Q[67]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF808F808FFFFF808)) 
    \Q[67]_i_11__0 
       (.I0(\Q[31]_i_11__0_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[31]_i_14__0_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[17]_i_10__0_n_0 ),
        .I5(\Q[21]_i_10__0_n_0 ),
        .O(\Q[67]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFCFFFCAA)) 
    \Q[67]_i_12 
       (.I0(ALU_DIN1[23]),
        .I1(\custom_alu/int2fp/INT_VAL0 [23]),
        .I2(\custom_alu/int2fp/INT_VAL0 [22]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(ALU_DIN1[22]),
        .I5(\Q[29]_i_10_n_0 ),
        .O(\Q[67]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00070000)) 
    \Q[67]_i_12__0 
       (.I0(\Q[4]_i_13_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[67]_i_13__0_n_0 ),
        .I3(\Q[23]_i_13_n_0 ),
        .I4(\custom_alu/fp32_add/significand_sub_complement1 ),
        .O(\Q[67]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[67]_i_13 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[31]_i_11__0_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[31]_i_14__0_n_0 ),
        .O(\Q[67]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000015155550151)) 
    \Q[67]_i_13__0 
       (.I0(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I1(\Q[67]_i_14_n_0 ),
        .I2(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I3(\Q[8]_i_18_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I5(\Q[4]_i_15_n_0 ),
        .O(\Q[67]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[67]_i_14 
       (.I0(ALU_DIN2[8]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[8]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[4]_i_23_n_0 ),
        .O(\Q[67]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFB00FBFF0B000B)) 
    \Q[67]_i_14__0 
       (.I0(\Q[28]_i_18_n_0 ),
        .I1(\Q[17]_i_10__0_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[28]_i_11_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[17]_i_11__0_n_0 ),
        .O(\Q[67]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'hCC88CC88CF8ACC8A)) 
    \Q[67]_i_15 
       (.I0(\Q[67]_i_17_n_0 ),
        .I1(\Q[67]_i_18_n_0 ),
        .I2(\Q[26]_i_23_n_0 ),
        .I3(\Q[35]_i_20_n_0 ),
        .I4(\Q[35]_i_22_n_0 ),
        .I5(\Q[35]_i_24_n_0 ),
        .O(\Q[67]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h22222222AAAA2AAA)) 
    \Q[67]_i_16 
       (.I0(\Q[67]_i_19_n_0 ),
        .I1(\Q[69]_i_22_n_0 ),
        .I2(ALU_DIN1[0]),
        .I3(\Q[29]_i_18__0_n_0 ),
        .I4(\Q[67]_i_20_n_0 ),
        .I5(\Q[67]_i_21_n_0 ),
        .O(\Q[67]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FBEAEAEA)) 
    \Q[67]_i_17 
       (.I0(\Q[35]_i_24_n_0 ),
        .I1(\Q[35]_i_19_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[35]_i_21_n_0 ),
        .I5(\Q[17]_i_14_n_0 ),
        .O(\Q[67]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFEBAEEAA)) 
    \Q[67]_i_18 
       (.I0(\Q[17]_i_14_n_0 ),
        .I1(\Q[17]_i_11__0_n_0 ),
        .I2(\Q[28]_i_18_n_0 ),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[35]_i_21_n_0 ),
        .O(\Q[67]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4447474774777777)) 
    \Q[67]_i_19 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_22_n_0 ),
        .I2(\Q[35]_i_27_n_0 ),
        .I3(\Q[17]_i_15_n_0 ),
        .I4(\Q[35]_i_26_n_0 ),
        .I5(\Q[35]_i_28_n_0 ),
        .O(\Q[67]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[67]_i_1__0 
       (.I0(\Q[67]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[20]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[20]),
        .I5(\Q[67]_i_4_n_0 ),
        .O(\Q[67]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[67]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[20]),
        .I2(CRF_RD1_IBUF[20]),
        .I3(RF_RD1_IBUF[20]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[67]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFCFFFFFFFCFAFA)) 
    \Q[67]_i_20 
       (.I0(ALU_DIN1[5]),
        .I1(\custom_alu/int2fp/INT_VAL0 [5]),
        .I2(\Q[35]_i_29_n_0 ),
        .I3(\custom_alu/int2fp/INT_VAL0 [4]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(ALU_DIN1[4]),
        .O(\Q[67]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[67]_i_21 
       (.I0(\Q[29]_i_18__0_n_0 ),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[35]_i_32_n_0 ),
        .I3(\Q[35]_i_28_n_0 ),
        .I4(\Q[17]_i_15_n_0 ),
        .I5(\Q[47]_i_9_n_0 ),
        .O(\Q[67]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBABA)) 
    \Q[67]_i_3 
       (.I0(\Q[25]_i_2_n_0 ),
        .I1(\Q[25]_i_3_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\Q[67]_i_5_n_0 ),
        .I4(\Q[67]_i_6_n_0 ),
        .O(CUSTOM_ALU_OUT[20]));
  LUT6 #(
    .INIT(64'hAAAAAAAA80AA8080)) 
    \Q[67]_i_4 
       (.I0(\Q[78]_i_4_n_0 ),
        .I1(\Q[36]_i_3__0_n_0 ),
        .I2(D_MEM_DOUT_IBUF[20]),
        .I3(MEM_D_MEM_ALU_FINAL1),
        .I4(EX_MEM_Q[25]),
        .I5(\Q[36]_i_2__1_n_0 ),
        .O(\Q[67]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h02A20000FEAE0000)) 
    \Q[67]_i_5 
       (.I0(\custom_alu/fp2int/p_0_in [20]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [20]),
        .O(\Q[67]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFBBBBAAAAAAAA)) 
    \Q[67]_i_6 
       (.I0(EX_CUSTOM_ALU_SEL[27]),
        .I1(\Q[67]_i_7_n_0 ),
        .I2(\Q[67]_i_8_n_0 ),
        .I3(\Q[67]_i_9__0_n_0 ),
        .I4(\Q[26]_i_7_n_0 ),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[67]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000553FFFFF553F)) 
    \Q[67]_i_7 
       (.I0(\Q[28]_i_12_n_0 ),
        .I1(\Q[23]_i_13__0_n_0 ),
        .I2(\Q[35]_i_16_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[67]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8AAA8A8A8A8)) 
    \Q[67]_i_8 
       (.I0(\Q[67]_i_10__0_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[29]_i_7_n_0 ),
        .I3(\Q[67]_i_11__0_n_0 ),
        .I4(\Q[67]_i_12_n_0 ),
        .I5(\Q[67]_i_13_n_0 ),
        .O(\Q[67]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h0000656A)) 
    \Q[67]_i_8__0 
       (.I0(PSUM3__0_carry__0_i_10__2_n_0),
        .I1(ID_EX_Q[110]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(EX_RF_RD2[31]),
        .I4(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/significand_sub_complement1 ));
  LUT5 #(
    .INIT(32'h8AAA8A88)) 
    \Q[67]_i_9 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[8]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[4]_i_11_n_0 ),
        .O(\Q[67]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h008A008A00FF008A)) 
    \Q[67]_i_9__0 
       (.I0(\Q[67]_i_14__0_n_0 ),
        .I1(\Q[67]_i_15_n_0 ),
        .I2(\Q[22]_i_7__0_n_0 ),
        .I3(\Q[27]_i_13_n_0 ),
        .I4(\Q[69]_i_20_n_0 ),
        .I5(\Q[67]_i_16_n_0 ),
        .O(\Q[67]_i_9__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[68]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [4]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [68]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[68]_i_1__0 
       (.I0(\Q[68]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[21]),
        .I4(data1[21]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[68]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[68]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[21]),
        .I3(CRF_RD1_IBUF[21]),
        .I4(CRF_WD_OBUF[21]),
        .O(\Q[68]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[69]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [5]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [69]));
  LUT5 #(
    .INIT(32'h44440400)) 
    \Q[69]_i_10 
       (.I0(\Q[27]_i_13_n_0 ),
        .I1(\Q[69]_i_20_n_0 ),
        .I2(\Q[69]_i_21_n_0 ),
        .I3(\Q[69]_i_22_n_0 ),
        .I4(\Q[69]_i_23_n_0 ),
        .O(\Q[69]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00F0FF0000DD)) 
    \Q[69]_i_11 
       (.I0(\Q[69]_i_24_n_0 ),
        .I1(\Q[69]_i_25_n_0 ),
        .I2(\Q[29]_i_10_n_0 ),
        .I3(\Q[35]_i_17_n_0 ),
        .I4(\Q[28]_i_12_n_0 ),
        .I5(\Q[23]_i_13__0_n_0 ),
        .O(\Q[69]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00FF474700FF47FF)) 
    \Q[69]_i_12 
       (.I0(\custom_alu/int2fp/INT_VAL0 [28]),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN1[28]),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[69]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \Q[69]_i_13 
       (.I0(\Q[69]_i_26_n_0 ),
        .I1(\Q[69]_i_27_n_0 ),
        .I2(\Q[69]_i_28_n_0 ),
        .I3(\Q[69]_i_29_n_0 ),
        .I4(\Q[69]_i_30_n_0 ),
        .I5(\Q[69]_i_31_n_0 ),
        .O(\Q[69]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40000000)) 
    \Q[69]_i_14 
       (.I0(\Q[69]_i_32_n_0 ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[30] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[23] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[29] ),
        .I4(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[24] ),
        .I5(\Q[69]_i_33_n_0 ),
        .O(\Q[69]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \Q[69]_i_15 
       (.I0(ALU_DIN1[18]),
        .I1(\custom_alu/int2fp/INT_VAL0 [18]),
        .I2(ALU_DIN1[16]),
        .I3(PSUM3__0_carry__0_i_10__2_n_0),
        .I4(\custom_alu/int2fp/INT_VAL0 [16]),
        .O(\Q[69]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBABF8A8FBAB08A80)) 
    \Q[69]_i_16 
       (.I0(\custom_alu/int2fp/INT_VAL0 [17]),
        .I1(ID_EX_Q[157]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__2_n_0 ),
        .I3(EX_RF_RD1[31]),
        .I4(ID_EX_Q[143]),
        .I5(EX_RF_RD1[17]),
        .O(\Q[69]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \Q[69]_i_17 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(EX_RF_RD1[15]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[141]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [15]),
        .O(\Q[69]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FA08)) 
    \Q[69]_i_18 
       (.I0(\Q[35]_i_21_n_0 ),
        .I1(\Q[35]_i_22_n_0 ),
        .I2(\Q[35]_i_20_n_0 ),
        .I3(\Q[35]_i_19_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[35]_i_24_n_0 ),
        .O(\Q[69]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00FF474700FF47FF)) 
    \Q[69]_i_19 
       (.I0(\custom_alu/int2fp/INT_VAL0 [13]),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN1[13]),
        .I3(\Q[17]_i_11__0_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[35]_i_20_n_0 ),
        .O(\Q[69]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAEA)) 
    \Q[69]_i_1__0 
       (.I0(\Q[69]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(D_MEM_ADDR_OBUF[22]),
        .I3(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I4(CUSTOM_ALU_OUT[22]),
        .I5(\Q[69]_i_4_n_0 ),
        .O(\Q[69]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[69]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[22]),
        .I2(CRF_RD1_IBUF[22]),
        .I3(RF_RD1_IBUF[22]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[69]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \Q[69]_i_20 
       (.I0(\Q[69]_i_15_n_0 ),
        .I1(\Q[69]_i_16_n_0 ),
        .I2(\Q[35]_i_21_n_0 ),
        .I3(\Q[29]_i_19__0_n_0 ),
        .I4(\Q[17]_i_14_n_0 ),
        .I5(\Q[35]_i_24_n_0 ),
        .O(\Q[69]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h4757475746564657)) 
    \Q[69]_i_21 
       (.I0(\Q[35]_i_28_n_0 ),
        .I1(\Q[35]_i_29_n_0 ),
        .I2(\Q[17]_i_15_n_0 ),
        .I3(\Q[29]_i_18__0_n_0 ),
        .I4(\Q[47]_i_9_n_0 ),
        .I5(\Q[69]_i_34_n_0 ),
        .O(\Q[69]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000440347)) 
    \Q[69]_i_22 
       (.I0(\custom_alu/int2fp/INT_VAL0 [8]),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN1[8]),
        .I3(\custom_alu/int2fp/INT_VAL0 [7]),
        .I4(ALU_DIN1[7]),
        .I5(\Q[35]_i_22_n_0 ),
        .O(\Q[69]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFF00B8B8FF00B800)) 
    \Q[69]_i_23 
       (.I0(\custom_alu/int2fp/INT_VAL0 [7]),
        .I1(\Q[63]_i_1__1_n_0 ),
        .I2(ALU_DIN1[7]),
        .I3(\Q[35]_i_27_n_0 ),
        .I4(\Q[35]_i_22_n_0 ),
        .I5(\Q[35]_i_29_n_0 ),
        .O(\Q[69]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h11DF111111DFDFDF)) 
    \Q[69]_i_24 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(\Q[29]_i_10_n_0 ),
        .I2(\Q[31]_i_14__0_n_0 ),
        .I3(\custom_alu/int2fp/INT_VAL0 [23]),
        .I4(\Q[63]_i_1__1_n_0 ),
        .I5(ALU_DIN1[23]),
        .O(\Q[69]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h000C000C000E0000)) 
    \Q[69]_i_25 
       (.I0(\Q[28]_i_11_n_0 ),
        .I1(\Q[31]_i_11__0_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[28]_i_13_n_0 ),
        .I4(\Q[31]_i_10__0_n_0 ),
        .I5(\Q[31]_i_14__0_n_0 ),
        .O(\Q[69]_i_25_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \Q[69]_i_26 
       (.I0(\custom_alu/fp32_mult/product_mantissa [9]),
        .I1(\custom_alu/fp32_mult/product_mantissa [8]),
        .I2(\custom_alu/fp32_mult/product_mantissa [11]),
        .I3(\custom_alu/fp32_mult/product_mantissa [10]),
        .O(\Q[69]_i_26_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \Q[69]_i_27 
       (.I0(\custom_alu/fp32_mult/product_mantissa [13]),
        .I1(\custom_alu/fp32_mult/product_mantissa [12]),
        .I2(\custom_alu/fp32_mult/product_mantissa [15]),
        .I3(\custom_alu/fp32_mult/product_mantissa [14]),
        .O(\Q[69]_i_27_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \Q[69]_i_28 
       (.I0(\custom_alu/fp32_mult/product_mantissa [1]),
        .I1(\custom_alu/fp32_mult/product_mantissa [0]),
        .I2(\custom_alu/fp32_mult/product_mantissa [3]),
        .I3(\custom_alu/fp32_mult/product_mantissa [2]),
        .O(\Q[69]_i_28_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \Q[69]_i_29 
       (.I0(\custom_alu/fp32_mult/product_mantissa [5]),
        .I1(\custom_alu/fp32_mult/product_mantissa [4]),
        .I2(\custom_alu/fp32_mult/product_mantissa [7]),
        .I3(\custom_alu/fp32_mult/product_mantissa [6]),
        .O(\Q[69]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAFBAAAAAAAA)) 
    \Q[69]_i_3 
       (.I0(\Q[27]_i_2__0_n_0 ),
        .I1(\Q[69]_i_5_n_0 ),
        .I2(\Q[69]_i_6_n_0 ),
        .I3(EX_CUSTOM_ALU_SEL[28]),
        .I4(\Q[69]_i_7_n_0 ),
        .I5(\Q[34]_i_5_n_0 ),
        .O(CUSTOM_ALU_OUT[22]));
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \Q[69]_i_30 
       (.I0(\custom_alu/fp32_mult/product_mantissa [21]),
        .I1(\custom_alu/fp32_mult/product_mantissa [22]),
        .I2(\custom_alu/fp32_mult/product_mantissa [20]),
        .O(\Q[69]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \Q[69]_i_31 
       (.I0(\custom_alu/fp32_mult/product_mantissa [17]),
        .I1(\custom_alu/fp32_mult/product_mantissa [16]),
        .I2(\custom_alu/fp32_mult/product_mantissa [19]),
        .I3(\custom_alu/fp32_mult/product_mantissa [18]),
        .O(\Q[69]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \Q[69]_i_32 
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[28] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[25] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[27] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[26] ),
        .O(\Q[69]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \Q[69]_i_33 
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[60] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[61] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[56] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[57] ),
        .I4(\Q[69]_i_35_n_0 ),
        .O(\Q[69]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h3055300033553355)) 
    \Q[69]_i_34 
       (.I0(ALU_DIN1[2]),
        .I1(\custom_alu/int2fp/INT_VAL0 [2]),
        .I2(\custom_alu/int2fp/INT_VAL0 [3]),
        .I3(\Q[63]_i_1__1_n_0 ),
        .I4(ALU_DIN1[3]),
        .I5(ALU_DIN1[0]),
        .O(\Q[69]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \Q[69]_i_35 
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[55] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[58] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[62] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[59] ),
        .O(\Q[69]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \Q[69]_i_4 
       (.I0(DIN1_FORWARD[0]),
        .I1(DIN1_FORWARD[1]),
        .I2(data1[22]),
        .O(\Q[69]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h02A2FFFFFEAEFFFF)) 
    \Q[69]_i_5 
       (.I0(\custom_alu/fp2int/p_0_in [22]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [22]),
        .O(\Q[69]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAA80000AAAAAAAA)) 
    \Q[69]_i_6 
       (.I0(\Q[27]_i_7_n_0 ),
        .I1(\Q[69]_i_9_n_0 ),
        .I2(\Q[69]_i_10_n_0 ),
        .I3(\Q[69]_i_11_n_0 ),
        .I4(\Q[26]_i_7_n_0 ),
        .I5(\Q[69]_i_12_n_0 ),
        .O(\Q[69]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \Q[69]_i_7 
       (.I0(\Q[69]_i_13_n_0 ),
        .I1(\Q[69]_i_14_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[28]),
        .I3(\custom_alu/fp32_mult/product_mantissa [22]),
        .I4(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .O(\Q[69]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAAAABFBFFFF)) 
    \Q[69]_i_8 
       (.I0(INT0_carry__4_i_4_n_0),
        .I1(EX_RF_RD1[22]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[148]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN1[23]),
        .O(\custom_alu/fp2int/p_0_in [22]));
  LUT6 #(
    .INIT(64'h4145404441454145)) 
    \Q[69]_i_9 
       (.I0(\Q[27]_i_13_n_0 ),
        .I1(\Q[69]_i_15_n_0 ),
        .I2(\Q[69]_i_16_n_0 ),
        .I3(\Q[69]_i_17_n_0 ),
        .I4(\Q[69]_i_18_n_0 ),
        .I5(\Q[69]_i_19_n_0 ),
        .O(\Q[69]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[6]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [6]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [5]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [6]));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[6]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[7] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/data23 [6]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\Q[6]_i_2_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [6]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[6]_i_1__1 
       (.I0(CUSTOM_ALU_OUT[1]),
        .I1(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I2(D_MEM_ADDR_OBUF[1]),
        .O(data0[1]));
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \Q[6]_i_1__2 
       (.I0(\Q[6]_i_2__0_n_0 ),
        .I1(\Q[11]_i_3__0_n_0 ),
        .I2(\Q[6]_i_3_n_0 ),
        .I3(\Q[11]_i_5__1_n_0 ),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(EX_MEM_Q[6]),
        .O(data1[1]));
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'h12)) 
    \Q[6]_i_1__3 
       (.I0(\Q[9]_i_4__1_n_0 ),
        .I1(STALL_COUNTER_D1),
        .I2(STALL_COUNTER_Q[6]),
        .O(STALL_COUNTER_D[6]));
  LUT5 #(
    .INIT(32'hBBB8B8B8)) 
    \Q[6]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\Q[6]_i_3__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [5]),
        .O(\Q[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[6]_i_2__0 
       (.I0(D_MEM_DOUT_IBUF[9]),
        .I1(D_MEM_DOUT_IBUF[1]),
        .I2(D_MEM_DOUT_IBUF[25]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[17]),
        .O(\Q[6]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[6]_i_3 
       (.I0(D_MEM_DOUT_IBUF[1]),
        .I1(D_MEM_DOUT_IBUF[17]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[25]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[9]),
        .O(\Q[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5555510100005101)) 
    \Q[6]_i_3__0 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .I1(\Q[6]_i_4_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [3]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [4]),
        .O(\Q[6]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h4444477777774777)) 
    \Q[6]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [17]),
        .I3(\custom_alu/fp32_add/sel0 [0]),
        .I4(\custom_alu/fp32_add/sel0 [18]),
        .I5(\custom_alu/fp32_add/sel0 [1]),
        .O(\Q[6]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[70]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [6]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [70]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[70]_i_1__0 
       (.I0(\Q[70]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(data0[23]),
        .I3(data1[23]),
        .I4(\Q[78]_i_4_n_0 ),
        .O(\Q[70]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[70]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[23]),
        .I2(CRF_RD1_IBUF[23]),
        .I3(RF_RD1_IBUF[23]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[70]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[71]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [7]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [71]));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[71]_i_10 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [5]),
        .O(\Q[71]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[71]_i_11 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [4]),
        .O(\Q[71]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[71]_i_1__0 
       (.I0(\Q[71]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[24]),
        .I4(data1[24]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[71]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[71]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[24]),
        .I3(CRF_RD1_IBUF[24]),
        .I4(CRF_WD_OBUF[24]),
        .O(\Q[71]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[71]_i_8 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [7]),
        .O(\Q[71]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[71]_i_9 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [6]),
        .O(\Q[71]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[72]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [8]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [72]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[72]_i_1__0 
       (.I0(\Q[72]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[25]),
        .I4(data1[25]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[72]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[72]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[25]),
        .I3(CRF_RD1_IBUF[25]),
        .I4(CRF_WD_OBUF[25]),
        .O(\Q[72]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[73]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [9]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [73]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[73]_i_1__0 
       (.I0(\Q[73]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(data0[26]),
        .I3(data1[26]),
        .I4(\Q[78]_i_4_n_0 ),
        .O(\Q[73]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[73]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[26]),
        .I2(CRF_RD1_IBUF[26]),
        .I3(RF_RD1_IBUF[26]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[73]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[74]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [10]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [74]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[74]_i_1__0 
       (.I0(\Q[74]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[27]),
        .I4(data1[27]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[74]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[74]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[27]),
        .I3(CRF_RD1_IBUF[27]),
        .I4(CRF_WD_OBUF[27]),
        .O(\Q[74]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[75]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [11]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [75]));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[75]_i_10 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [9]),
        .O(\Q[75]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[75]_i_11 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [8]),
        .O(\Q[75]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[75]_i_1__0 
       (.I0(\Q[75]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[28]),
        .I4(data1[28]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[75]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[75]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[28]),
        .I3(CRF_RD1_IBUF[28]),
        .I4(CRF_WD_OBUF[28]),
        .O(\Q[75]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[75]_i_8 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [11]),
        .O(\Q[75]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[75]_i_9 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [10]),
        .O(\Q[75]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[76]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [12]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [76]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[76]_i_1__0 
       (.I0(\Q[76]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[29]),
        .I4(data1[29]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[76]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[76]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[29]),
        .I3(CRF_RD1_IBUF[29]),
        .I4(CRF_WD_OBUF[29]),
        .O(\Q[76]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[77]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [13]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [77]));
  LUT6 #(
    .INIT(64'hFFFFF111F111F111)) 
    \Q[77]_i_1__0 
       (.I0(\Q[77]_i_2_n_0 ),
        .I1(\Q[77]_i_3_n_0 ),
        .I2(\Q[78]_i_3_n_0 ),
        .I3(data0[30]),
        .I4(data1[30]),
        .I5(\Q[78]_i_4_n_0 ),
        .O(\Q[77]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'h0123CDEF)) 
    \Q[77]_i_2 
       (.I0(CUSTOM_RS1),
        .I1(DIN1_FORWARD[2]),
        .I2(RF_RD1_IBUF[30]),
        .I3(CRF_RD1_IBUF[30]),
        .I4(CRF_WD_OBUF[30]),
        .O(\Q[77]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01000001)) 
    \Q[77]_i_3 
       (.I0(\Q[77]_i_4_n_0 ),
        .I1(\Q[77]_i_5_n_0 ),
        .I2(\Q[77]_i_6_n_0 ),
        .I3(EX_MEM_Q[0]),
        .I4(CRF_RA1_OBUF[0]),
        .I5(DIN1_FORWARD[0]),
        .O(\Q[77]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \Q[77]_i_4 
       (.I0(CRF_RA1_OBUF[3]),
        .I1(EX_MEM_Q[3]),
        .I2(CRF_RA1_OBUF[1]),
        .I3(EX_MEM_Q[1]),
        .I4(EX_MEM_Q[4]),
        .I5(CRF_RA1_OBUF[4]),
        .O(\Q[77]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT4 #(
    .INIT(16'h6FF6)) 
    \Q[77]_i_5 
       (.I0(CUSTOM_RS1),
        .I1(MEM_CUSTOM_RD),
        .I2(CRF_RA1_OBUF[2]),
        .I3(EX_MEM_Q[2]),
        .O(\Q[77]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \Q[77]_i_6 
       (.I0(EX_MEM_Q[3]),
        .I1(EX_MEM_Q[4]),
        .I2(EX_MEM_Q[2]),
        .I3(EX_MEM_Q[1]),
        .I4(EX_MEM_Q[0]),
        .I5(EX_MEM_Q[38]),
        .O(\Q[77]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[78]_i_1 
       (.I0(\custom_alu/fp32_add/significand_sub0 [14]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [78]));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT5 #(
    .INIT(32'hFFFF6FF6)) 
    \Q[78]_i_10 
       (.I0(EX_MEM_Q[2]),
        .I1(CRF_RA1_OBUF[2]),
        .I2(MEM_CUSTOM_RD),
        .I3(CUSTOM_RS1),
        .I4(\Q[78]_i_16_n_0 ),
        .O(\Q[78]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \Q[78]_i_11 
       (.I0(CRF_RA1_OBUF[4]),
        .I1(CRF_WA_OBUF[4]),
        .I2(CRF_RA1_OBUF[3]),
        .I3(CRF_WA_OBUF[3]),
        .I4(CRF_WA_OBUF[2]),
        .I5(CRF_RA1_OBUF[2]),
        .O(\Q[78]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hBEFFFFBE)) 
    \Q[78]_i_12 
       (.I0(\Q[78]_i_17_n_0 ),
        .I1(CRF_RA1_OBUF[4]),
        .I2(ID_EX_Q[4]),
        .I3(ID_EX_Q[0]),
        .I4(CRF_RA1_OBUF[0]),
        .O(\Q[78]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h6FF6)) 
    \Q[78]_i_13 
       (.I0(ID_EX_Q[1]),
        .I1(CRF_RA1_OBUF[1]),
        .I2(ID_EX_Q[3]),
        .I3(CRF_RA1_OBUF[3]),
        .O(\Q[78]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h6FF6)) 
    \Q[78]_i_14 
       (.I0(CRF_RA1_OBUF[0]),
        .I1(CRF_WA_OBUF[0]),
        .I2(CRF_RA1_OBUF[1]),
        .I3(CRF_WA_OBUF[1]),
        .O(\Q[78]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \Q[78]_i_15 
       (.I0(CRF_WA_OBUF[3]),
        .I1(CRF_WA_OBUF[4]),
        .I2(CRF_WA_OBUF[2]),
        .I3(CRF_WA_OBUF[1]),
        .I4(CRF_WA_OBUF[0]),
        .I5(MEM_WB_Q),
        .O(\Q[78]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hF6)) 
    \Q[78]_i_16 
       (.I0(CRF_RA1_OBUF[0]),
        .I1(EX_MEM_Q[0]),
        .I2(\Q[77]_i_6_n_0 ),
        .O(\Q[78]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \Q[78]_i_17 
       (.I0(ID_EX_Q[3]),
        .I1(ID_EX_Q[4]),
        .I2(ID_EX_Q[2]),
        .I3(ID_EX_Q[1]),
        .I4(ID_EX_Q[0]),
        .I5(ID_EX_Q[113]),
        .O(\Q[78]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \Q[78]_i_1__0 
       (.I0(\Q[78]_i_2_n_0 ),
        .I1(\Q[78]_i_3_n_0 ),
        .I2(data0[31]),
        .I3(data1[31]),
        .I4(\Q[78]_i_4_n_0 ),
        .O(\Q[78]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D8D8DD88)) 
    \Q[78]_i_2 
       (.I0(DIN1_FORWARD[2]),
        .I1(CRF_WD_OBUF[31]),
        .I2(CRF_RD1_IBUF[31]),
        .I3(RF_RD1_IBUF[31]),
        .I4(CUSTOM_RS1),
        .I5(\Q[77]_i_3_n_0 ),
        .O(\Q[78]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \Q[78]_i_3 
       (.I0(\Q[77]_i_3_n_0 ),
        .I1(DIN1_FORWARD[0]),
        .O(\Q[78]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[78]_i_4 
       (.I0(DIN1_FORWARD[1]),
        .I1(DIN1_FORWARD[0]),
        .O(\Q[78]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00005554)) 
    \Q[78]_i_5 
       (.I0(\Q[78]_i_9_n_0 ),
        .I1(\Q[78]_i_10_n_0 ),
        .I2(DIN1_FORWARD[0]),
        .I3(\Q[77]_i_4_n_0 ),
        .I4(\Q[78]_i_11_n_0 ),
        .O(DIN1_FORWARD[2]));
  LUT3 #(
    .INIT(8'hF4)) 
    \Q[78]_i_6 
       (.I0(I_MEM_DOUT_IBUF[28]),
        .I1(\Q[27]_i_2_n_0 ),
        .I2(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .O(CUSTOM_RS1));
  LUT6 #(
    .INIT(64'h1001000000001001)) 
    \Q[78]_i_7 
       (.I0(\Q[78]_i_12_n_0 ),
        .I1(\Q[78]_i_13_n_0 ),
        .I2(ID_EX_Q[2]),
        .I3(CRF_RA1_OBUF[2]),
        .I4(EX_CUSTOM_RD),
        .I5(CUSTOM_RS1),
        .O(DIN1_FORWARD[0]));
  LUT6 #(
    .INIT(64'h0000000000000009)) 
    \Q[78]_i_8 
       (.I0(CRF_RA1_OBUF[0]),
        .I1(EX_MEM_Q[0]),
        .I2(\Q[77]_i_6_n_0 ),
        .I3(\Q[77]_i_5_n_0 ),
        .I4(DIN1_FORWARD[0]),
        .I5(\Q[77]_i_4_n_0 ),
        .O(DIN1_FORWARD[1]));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT4 #(
    .INIT(16'hEFFE)) 
    \Q[78]_i_9 
       (.I0(\Q[78]_i_14_n_0 ),
        .I1(\Q[78]_i_15_n_0 ),
        .I2(WB_CUSTOM_RD),
        .I3(CUSTOM_RS1),
        .O(\Q[78]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEAAAEAAAEAAA)) 
    \Q[79]_i_1 
       (.I0(\Q[79]_i_2_n_0 ),
        .I1(I_MEM_DOUT_FILTERED[7]),
        .I2(\Q[79]_i_3_n_0 ),
        .I3(\Q[112]_i_2_n_0 ),
        .I4(CRF_RA2_OBUF[0]),
        .I5(\Q[79]_i_4_n_0 ),
        .O(ID_IMMEDIATE[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[79]_i_10 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [13]),
        .O(\Q[79]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[79]_i_11 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [12]),
        .O(\Q[79]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[79]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [15]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [79]));
  LUT6 #(
    .INIT(64'h8AAA8AAAA280A080)) 
    \Q[79]_i_2 
       (.I0(CRF_RA2_OBUF[0]),
        .I1(I_MEM_DOUT_FILTERED[4]),
        .I2(I_MEM_DOUT_FILTERED[6]),
        .I3(I_MEM_DOUT_FILTERED[2]),
        .I4(\Q[160]_i_2_n_0 ),
        .I5(I_MEM_DOUT_FILTERED[3]),
        .O(\Q[79]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    \Q[79]_i_3 
       (.I0(I_MEM_DOUT_IBUF[5]),
        .I1(I_MEM_DOUT_IBUF[4]),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[3]),
        .O(\Q[79]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT4 #(
    .INIT(16'hCDFD)) 
    \Q[79]_i_4 
       (.I0(I_MEM_DOUT_IBUF[5]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[4]),
        .I3(I_MEM_DOUT_IBUF[2]),
        .O(\Q[79]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[79]_i_8 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [15]),
        .O(\Q[79]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[79]_i_9 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [14]),
        .O(\Q[79]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[7]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [7]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [6]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [7]));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[7]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[8] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\Q[7]_i_2_n_0 ),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [7]));
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[7]_i_1__1 
       (.I0(CUSTOM_ALU_OUT[2]),
        .I1(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I2(D_MEM_ADDR_OBUF[2]),
        .O(data0[2]));
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \Q[7]_i_1__2 
       (.I0(\Q[7]_i_2__0_n_0 ),
        .I1(\Q[11]_i_3__0_n_0 ),
        .I2(\Q[7]_i_3__0_n_0 ),
        .I3(\Q[11]_i_5__1_n_0 ),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(EX_MEM_Q[7]),
        .O(data1[2]));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT4 #(
    .INIT(16'h0708)) 
    \Q[7]_i_1__3 
       (.I0(STALL_COUNTER_Q[6]),
        .I1(\Q[9]_i_4__1_n_0 ),
        .I2(STALL_COUNTER_D1),
        .I3(STALL_COUNTER_Q[7]),
        .O(STALL_COUNTER_D[7]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[7]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\Q[7]_i_3_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\custom_alu/fp32_add/data23 [7]),
        .O(\Q[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[7]_i_2__0 
       (.I0(D_MEM_DOUT_IBUF[10]),
        .I1(D_MEM_DOUT_IBUF[2]),
        .I2(D_MEM_DOUT_IBUF[26]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[18]),
        .O(\Q[7]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'hFF8B008B)) 
    \Q[7]_i_3 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .I1(\custom_alu/fp32_add/sel0 [21]),
        .I2(\Q[7]_i_4_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [6]),
        .O(\Q[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[7]_i_3__0 
       (.I0(D_MEM_DOUT_IBUF[2]),
        .I1(D_MEM_DOUT_IBUF[18]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[26]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[10]),
        .O(\Q[7]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h47444777)) 
    \Q[7]_i_4 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [20]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [19]),
        .I4(\Q[7]_i_5_n_0 ),
        .O(\Q[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[7]_i_5 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [17]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [16]),
        .O(\Q[7]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT5 #(
    .INIT(32'hFF202020)) 
    \Q[80]_i_1 
       (.I0(I_MEM_DOUT_IBUF[8]),
        .I1(EX_BR_TAKEN),
        .I2(\Q[83]_i_2_n_0 ),
        .I3(CRF_RA2_OBUF[1]),
        .I4(\Q[83]_i_3_n_0 ),
        .O(ID_IMMEDIATE[1]));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[80]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [16]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [80]));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'hFF202020)) 
    \Q[81]_i_1 
       (.I0(I_MEM_DOUT_IBUF[9]),
        .I1(EX_BR_TAKEN),
        .I2(\Q[83]_i_2_n_0 ),
        .I3(CRF_RA2_OBUF[2]),
        .I4(\Q[83]_i_3_n_0 ),
        .O(ID_IMMEDIATE[2]));
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[81]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [17]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [81]));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT5 #(
    .INIT(32'hFF202020)) 
    \Q[82]_i_1 
       (.I0(I_MEM_DOUT_IBUF[10]),
        .I1(EX_BR_TAKEN),
        .I2(\Q[83]_i_2_n_0 ),
        .I3(CRF_RA2_OBUF[3]),
        .I4(\Q[83]_i_3_n_0 ),
        .O(ID_IMMEDIATE[3]));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[82]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [18]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [82]));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT5 #(
    .INIT(32'hFF202020)) 
    \Q[83]_i_1 
       (.I0(I_MEM_DOUT_IBUF[11]),
        .I1(EX_BR_TAKEN),
        .I2(\Q[83]_i_2_n_0 ),
        .I3(CRF_RA2_OBUF[4]),
        .I4(\Q[83]_i_3_n_0 ),
        .O(ID_IMMEDIATE[4]));
  LUT5 #(
    .INIT(32'h8A888AAA)) 
    \Q[83]_i_10 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[20]_i_12__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_13__1_n_0 ),
        .O(\Q[83]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h8A888AAA)) 
    \Q[83]_i_11 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[20]_i_13__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_14__1_n_0 ),
        .O(\Q[83]_i_11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[83]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [19]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [83]));
  LUT6 #(
    .INIT(64'h00000000CDCDCDCF)) 
    \Q[83]_i_2 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[3]),
        .I3(\Q[160]_i_2_n_0 ),
        .I4(I_MEM_DOUT_IBUF[6]),
        .I5(\Q[161]_i_4_n_0 ),
        .O(\Q[83]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF5FFF5FFFFF7F7F7)) 
    \Q[83]_i_3 
       (.I0(\Q[125]_i_2_n_0 ),
        .I1(I_MEM_DOUT_FILTERED[5]),
        .I2(I_MEM_DOUT_FILTERED[3]),
        .I3(I_MEM_DOUT_FILTERED[2]),
        .I4(\Q[160]_i_2_n_0 ),
        .I5(I_MEM_DOUT_FILTERED[4]),
        .O(\Q[83]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h8A888AAA)) 
    \Q[83]_i_8 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[23]_i_15_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_11__1_n_0 ),
        .O(\Q[83]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h8A888AAA)) 
    \Q[83]_i_9 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[20]_i_11__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_12__1_n_0 ),
        .O(\Q[83]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[84]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[25]),
        .O(ID_IMMEDIATE[5]));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[84]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [20]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [84]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[85]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[26]),
        .O(ID_IMMEDIATE[6]));
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[85]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [21]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [85]));
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[86]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[27]),
        .O(ID_IMMEDIATE[7]));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[86]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [22]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [86]));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[87]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[28]),
        .O(ID_IMMEDIATE[8]));
  LUT6 #(
    .INIT(64'hAA8A8888AA8AAAAA)) 
    \Q[87]_i_10 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[23]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I5(\Q[23]_i_14_n_0 ),
        .O(\Q[87]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h8A888AAA)) 
    \Q[87]_i_11 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[23]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[23]_i_15_n_0 ),
        .O(\Q[87]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFB8)) 
    \Q[87]_i_12 
       (.I0(ALU_DIN2[30]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[30]),
        .I3(\custom_alu/fp32_add/p_0_in [4]),
        .I4(\custom_alu/fp32_add/p_0_in [6]),
        .I5(\custom_alu/fp32_add/p_0_in [5]),
        .O(\Q[87]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[87]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [23]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [87]));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFE)) 
    \Q[87]_i_4 
       (.I0(\Q[87]_i_12_n_0 ),
        .I1(\custom_alu/fp32_add/p_0_in [2]),
        .I2(\custom_alu/fp32_add/p_0_in [3]),
        .I3(\custom_alu/fp32_add/p_0_in [1]),
        .I4(\custom_alu/fp32_add/p_0_in [0]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [23]),
        .O(\Q[87]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[87]_i_8 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [23]),
        .O(\Q[87]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[87]_i_9 
       (.I0(\custom_alu/fp32_add/significand_sub_complement1 ),
        .I1(\custom_alu/fp32_add/significand_b_add_sub [22]),
        .O(\Q[87]_i_9_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[88]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[29]),
        .O(ID_IMMEDIATE[9]));
  LUT2 #(
    .INIT(4'h2)) 
    \Q[88]_i_1__0 
       (.I0(\custom_alu/fp32_add/significand_sub0 [24]),
        .I1(\Q[88]_i_3_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [88]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF6FF6)) 
    \Q[88]_i_3 
       (.I0(\custom_alu/fp32_add/exp_b_add_sub [6]),
        .I1(\custom_alu/fp32_add/p_0_in [6]),
        .I2(\custom_alu/fp32_add/exp_b_add_sub [7]),
        .I3(\custom_alu/fp32_add/p_0_in [7]),
        .I4(\Q[88]_i_4_n_0 ),
        .I5(\Q[88]_i_5_n_0 ),
        .O(\Q[88]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \Q[88]_i_4 
       (.I0(\custom_alu/fp32_add/p_0_in [0]),
        .I1(\custom_alu/fp32_add/exp_b_add_sub [0]),
        .I2(\custom_alu/fp32_add/exp_b_add_sub [1]),
        .I3(\custom_alu/fp32_add/p_0_in [1]),
        .I4(\custom_alu/fp32_add/exp_b_add_sub [2]),
        .I5(\custom_alu/fp32_add/p_0_in [2]),
        .O(\Q[88]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \Q[88]_i_5 
       (.I0(\custom_alu/fp32_add/exp_b_add_sub [4]),
        .I1(\custom_alu/fp32_add/p_0_in [4]),
        .I2(\custom_alu/fp32_add/exp_b_add_sub [5]),
        .I3(\custom_alu/fp32_add/p_0_in [5]),
        .I4(\custom_alu/fp32_add/p_0_in [3]),
        .I5(\custom_alu/fp32_add/exp_b_add_sub [3]),
        .O(\Q[88]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \Q[89]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[30]),
        .O(ID_IMMEDIATE[10]));
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[8]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [8]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [7]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [8]));
  LUT6 #(
    .INIT(64'h4744477747774777)) 
    \Q[8]_i_10 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\custom_alu/fp32_add/sel0 [0]),
        .O(\Q[8]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h0000CCA0)) 
    \Q[8]_i_10__0 
       (.I0(ALU_DIN1[0]),
        .I1(\Q[47]_i_9_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[31]_i_14__0_n_0 ),
        .I4(\Q[31]_i_13__0_n_0 ),
        .O(\Q[8]_i_10__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[8]_i_11 
       (.I0(\Q[12]_i_15_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[8]_i_15_n_0 ),
        .O(\Q[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \Q[8]_i_12 
       (.I0(\Q[12]_i_18_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[12]_i_19_n_0 ),
        .I3(\Q[12]_i_16_n_0 ),
        .I4(\Q[8]_i_16_n_0 ),
        .I5(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[8]_i_12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \Q[8]_i_13 
       (.I0(\Q[12]_i_17_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[8]_i_17_n_0 ),
        .O(\Q[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \Q[8]_i_14 
       (.I0(\Q[12]_i_19_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [2]),
        .I2(\Q[8]_i_18_n_0 ),
        .I3(\Q[12]_i_16_n_0 ),
        .I4(\Q[8]_i_16_n_0 ),
        .I5(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(\Q[8]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[8]_i_15 
       (.I0(ALU_DIN2[15]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[15]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[8]_i_19_n_0 ),
        .O(\Q[8]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[8]_i_16 
       (.I0(ALU_DIN2[14]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[14]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[8]_i_20_n_0 ),
        .O(\Q[8]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[8]_i_17 
       (.I0(ALU_DIN2[13]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[13]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[8]_i_21_n_0 ),
        .O(\Q[8]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \Q[8]_i_18 
       (.I0(ALU_DIN2[12]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN1[12]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [3]),
        .I5(\Q[8]_i_22_n_0 ),
        .O(\Q[8]_i_18_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT5 #(
    .INIT(32'h00B8FFB8)) 
    \Q[8]_i_19 
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN2[7]),
        .I3(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I4(\Q[23]_i_22_n_0 ),
        .O(\Q[8]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[8]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[9] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\custom_alu/fp32_add/data23 [8]),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\Q[8]_i_3__0_n_0 ),
        .I5(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [8]));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[8]_i_1__1 
       (.I0(\Q[8]_i_2_n_0 ),
        .I1(\Q[8]_i_3__1_n_0 ),
        .I2(\Q[8]_i_4_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[3]),
        .O(data0[3]));
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \Q[8]_i_1__2 
       (.I0(\Q[8]_i_2__0_n_0 ),
        .I1(\Q[11]_i_3__0_n_0 ),
        .I2(\Q[8]_i_3__2_n_0 ),
        .I3(\Q[11]_i_5__1_n_0 ),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(EX_MEM_Q[8]),
        .O(data1[3]));
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT5 #(
    .INIT(32'h007F0080)) 
    \Q[8]_i_1__3 
       (.I0(STALL_COUNTER_Q[7]),
        .I1(\Q[9]_i_4__1_n_0 ),
        .I2(STALL_COUNTER_Q[6]),
        .I3(STALL_COUNTER_D1),
        .I4(STALL_COUNTER_Q[8]),
        .O(STALL_COUNTER_D[8]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[8]_i_2 
       (.I0(\custom_alu/MULT [3]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [35]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [3]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \Q[8]_i_20 
       (.I0(ALU_DIN1[22]),
        .I1(ALU_DIN2[22]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I3(ALU_DIN1[6]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[6]),
        .O(\Q[8]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \Q[8]_i_21 
       (.I0(ALU_DIN1[21]),
        .I1(ALU_DIN2[21]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I3(ALU_DIN1[5]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN2[5]),
        .O(\Q[8]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \Q[8]_i_22 
       (.I0(ALU_DIN1[20]),
        .I1(ALU_DIN2[20]),
        .I2(\custom_alu/fp32_add/p_1_in__0 [4]),
        .I3(ALU_DIN1[4]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(op_a2_carry_i_9_n_0),
        .O(\Q[8]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[8]_i_2__0 
       (.I0(D_MEM_DOUT_IBUF[11]),
        .I1(D_MEM_DOUT_IBUF[3]),
        .I2(D_MEM_DOUT_IBUF[27]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[19]),
        .O(\Q[8]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[8]_i_2__1 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[8]),
        .I2(STALL_EN),
        .I3(IF_PC2[8]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[8] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[8]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[8]_i_3 
       (.I0(\Q[8]_i_11_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\Q[12]_i_13_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[12]_i_14__0_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [7]));
  LUT5 #(
    .INIT(32'hBBB8B8B8)) 
    \Q[8]_i_3__0 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\Q[8]_i_8__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [7]),
        .O(\Q[8]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \Q[8]_i_3__1 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [3]),
        .O(\Q[8]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[8]_i_3__2 
       (.I0(D_MEM_DOUT_IBUF[3]),
        .I1(D_MEM_DOUT_IBUF[19]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[27]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[11]),
        .O(\Q[8]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[8]_i_3__3 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[7]),
        .I2(STALL_EN),
        .I3(IF_PC2[7]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[7] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[8]_i_3__3_n_0 ));
  LUT6 #(
    .INIT(64'h00FC00B8003000B8)) 
    \Q[8]_i_4 
       (.I0(INT0_carry_i_11_n_0),
        .I1(EX_CUSTOM_ALU_SEL[27]),
        .I2(\Q[8]_i_5__1_n_0 ),
        .I3(EX_CUSTOM_ALU_SEL[28]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/fp2int/INT0 [3]),
        .O(\Q[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[8]_i_4__0 
       (.I0(\Q[8]_i_12_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[8]_i_11_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[12]_i_13_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [6]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[8]_i_4__1 
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .O(\Q[8]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[8]_i_4__2 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[6]),
        .I2(STALL_EN),
        .I3(IF_PC2[6]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[6] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[8]_i_4__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \Q[8]_i_5 
       (.I0(\Q[8]_i_13_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I2(\Q[8]_i_11_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[8]_i_12_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [5]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[8]_i_5__0 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .O(\Q[8]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000A8080202AA0A)) 
    \Q[8]_i_5__1 
       (.I0(EX_CUSTOM_ALU_SEL[26]),
        .I1(\Q[26]_i_15__0_n_0 ),
        .I2(\Q[28]_i_6_n_0 ),
        .I3(\Q[35]_i_21_n_0 ),
        .I4(\Q[8]_i_6__1_n_0 ),
        .I5(\Q[8]_i_7__0_n_0 ),
        .O(\Q[8]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A808A8A8080)) 
    \Q[8]_i_5__2 
       (.I0(RSTn_IBUF),
        .I1(ID_PC[5]),
        .I2(STALL_EN),
        .I3(IF_PC2[5]),
        .I4(\FF_IF_ID_PCADD/Q_reg_n_0_[5] ),
        .I5(EX_BR_TAKEN),
        .O(\Q[8]_i_5__2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \Q[8]_i_6 
       (.I0(\Q[8]_i_14_n_0 ),
        .I1(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I2(\Q[8]_i_13_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\Q[8]_i_11_n_0 ),
        .I5(\Q[23]_i_13_n_0 ),
        .O(\custom_alu/fp32_add/significand_b_add_sub [4]));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[8]_i_6__0 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .O(\Q[8]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000777)) 
    \Q[8]_i_6__1 
       (.I0(\Q[28]_i_7_n_0 ),
        .I1(\Q[35]_i_27_n_0 ),
        .I2(\Q[35]_i_18_n_0 ),
        .I3(\Q[35]_i_22_n_0 ),
        .I4(\Q[28]_i_6_n_0 ),
        .O(\Q[8]_i_6__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[8]_i_7 
       (.I0(\custom_alu/fp32_add/sel0 [5]),
        .O(\Q[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h888A8A8A88888888)) 
    \Q[8]_i_7__0 
       (.I0(\Q[8]_i_8_n_0 ),
        .I1(\Q[8]_i_9__0_n_0 ),
        .I2(\Q[8]_i_10__0_n_0 ),
        .I3(\Q[35]_i_32_n_0 ),
        .I4(\Q[31]_i_13__0_n_0 ),
        .I5(\Q[29]_i_5__0_n_0 ),
        .O(\Q[8]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000535FFFFF535F)) 
    \Q[8]_i_8 
       (.I0(\Q[35]_i_29_n_0 ),
        .I1(\Q[35]_i_28_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[23]_i_13__0_n_0 ),
        .I4(\Q[35]_i_17_n_0 ),
        .I5(\Q[35]_i_26_n_0 ),
        .O(\Q[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5555510100005101)) 
    \Q[8]_i_8__0 
       (.I0(\custom_alu/fp32_add/sel0 [22]),
        .I1(\Q[8]_i_9_n_0 ),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [5]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [6]),
        .O(\Q[8]_i_8__0_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[8]_i_9 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [18]),
        .I4(\Q[8]_i_10_n_0 ),
        .O(\Q[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF02F2)) 
    \Q[8]_i_9__0 
       (.I0(\Q[28]_i_20_n_0 ),
        .I1(\Q[29]_i_18__0_n_0 ),
        .I2(\Q[29]_i_10_n_0 ),
        .I3(\Q[17]_i_15_n_0 ),
        .I4(\Q[29]_i_7_n_0 ),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[8]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEFEEEEE)) 
    \Q[90]_i_1 
       (.I0(\Q[90]_i_2_n_0 ),
        .I1(\Q[90]_i_3_n_0 ),
        .I2(\Q[90]_i_4_n_0 ),
        .I3(EX_BR_TAKEN),
        .I4(I_MEM_DOUT_IBUF[7]),
        .I5(\Q[90]_i_5_n_0 ),
        .O(ID_IMMEDIATE[11]));
  LUT6 #(
    .INIT(64'h00000000BA00AA00)) 
    \Q[90]_i_2 
       (.I0(\Q[90]_i_6_n_0 ),
        .I1(\Q[125]_i_2_n_0 ),
        .I2(CRF_RA2_OBUF[0]),
        .I3(I_MEM_DOUT_FILTERED[3]),
        .I4(I_MEM_DOUT_FILTERED[5]),
        .I5(I_MEM_DOUT_FILTERED[4]),
        .O(\Q[90]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h1111000033F30000)) 
    \Q[90]_i_3 
       (.I0(I_MEM_DOUT_FILTERED[5]),
        .I1(I_MEM_DOUT_FILTERED[4]),
        .I2(\Q[109]_i_3_n_0 ),
        .I3(I_MEM_DOUT_FILTERED[2]),
        .I4(I_MEM_DOUT_IBUF[31]),
        .I5(I_MEM_DOUT_FILTERED[6]),
        .O(\Q[90]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \Q[90]_i_4 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(I_MEM_DOUT_IBUF[4]),
        .I2(I_MEM_DOUT_IBUF[5]),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(EX_BR_TAKEN),
        .I5(I_MEM_DOUT_IBUF[6]),
        .O(\Q[90]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFAC000005A000000)) 
    \Q[90]_i_5 
       (.I0(I_MEM_DOUT_FILTERED[3]),
        .I1(\Q[109]_i_3_n_0 ),
        .I2(I_MEM_DOUT_FILTERED[6]),
        .I3(I_MEM_DOUT_FILTERED[2]),
        .I4(I_MEM_DOUT_IBUF[31]),
        .I5(I_MEM_DOUT_FILTERED[4]),
        .O(\Q[90]_i_5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \Q[90]_i_6 
       (.I0(I_MEM_DOUT_IBUF[31]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[2]),
        .O(\Q[90]_i_6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \Q[91]_i_1 
       (.I0(I_MEM_DOUT_IBUF[12]),
        .I1(\Q[98]_i_2_n_0 ),
        .I2(\Q[98]_i_3_n_0 ),
        .O(ID_IMMEDIATE[12]));
  LUT6 #(
    .INIT(64'hFFFFBAAABAAABAAA)) 
    \Q[92]_i_1 
       (.I0(\Q[92]_i_2_n_0 ),
        .I1(I_MEM_DOUT_FILTERED[2]),
        .I2(I_MEM_DOUT_IBUF[31]),
        .I3(I_MEM_DOUT_FILTERED[5]),
        .I4(I_MEM_DOUT_IBUF[13]),
        .I5(\Q[98]_i_2_n_0 ),
        .O(ID_IMMEDIATE[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFCCCC888C)) 
    \Q[92]_i_2 
       (.I0(\Q[98]_i_4_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(I_MEM_DOUT_IBUF[12]),
        .I3(I_MEM_DOUT_FILTERED[2]),
        .I4(I_MEM_DOUT_IBUF[13]),
        .I5(\Q[92]_i_3_n_0 ),
        .O(\Q[92]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT5 #(
    .INIT(32'h04080000)) 
    \Q[92]_i_3 
       (.I0(I_MEM_DOUT_IBUF[6]),
        .I1(I_MEM_DOUT_IBUF[2]),
        .I2(EX_BR_TAKEN),
        .I3(I_MEM_DOUT_IBUF[3]),
        .I4(I_MEM_DOUT_IBUF[31]),
        .O(\Q[92]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \Q[93]_i_1 
       (.I0(I_MEM_DOUT_IBUF[14]),
        .I1(\Q[98]_i_2_n_0 ),
        .I2(\Q[98]_i_3_n_0 ),
        .O(ID_IMMEDIATE[14]));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \Q[94]_i_1 
       (.I0(CRF_RA1_OBUF[0]),
        .I1(\Q[98]_i_2_n_0 ),
        .I2(\Q[98]_i_3_n_0 ),
        .O(ID_IMMEDIATE[15]));
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \Q[95]_i_1 
       (.I0(CRF_RA1_OBUF[1]),
        .I1(\Q[98]_i_2_n_0 ),
        .I2(\Q[98]_i_3_n_0 ),
        .O(ID_IMMEDIATE[16]));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \Q[96]_i_1 
       (.I0(CRF_RA1_OBUF[2]),
        .I1(\Q[98]_i_2_n_0 ),
        .I2(\Q[98]_i_3_n_0 ),
        .O(ID_IMMEDIATE[17]));
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \Q[97]_i_1 
       (.I0(CRF_RA1_OBUF[3]),
        .I1(\Q[98]_i_2_n_0 ),
        .I2(\Q[98]_i_3_n_0 ),
        .O(ID_IMMEDIATE[18]));
  LUT3 #(
    .INIT(8'hF8)) 
    \Q[98]_i_1 
       (.I0(CRF_RA1_OBUF[4]),
        .I1(\Q[98]_i_2_n_0 ),
        .I2(\Q[98]_i_3_n_0 ),
        .O(ID_IMMEDIATE[19]));
  LUT6 #(
    .INIT(64'h0003000008000000)) 
    \Q[98]_i_2 
       (.I0(I_MEM_DOUT_IBUF[5]),
        .I1(I_MEM_DOUT_IBUF[3]),
        .I2(EX_BR_TAKEN),
        .I3(I_MEM_DOUT_IBUF[6]),
        .I4(I_MEM_DOUT_IBUF[2]),
        .I5(I_MEM_DOUT_IBUF[4]),
        .O(\Q[98]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFEEFAEE00000000)) 
    \Q[98]_i_3 
       (.I0(\Q[98]_i_4_n_0 ),
        .I1(\Q[109]_i_3_n_0 ),
        .I2(I_MEM_DOUT_FILTERED[6]),
        .I3(I_MEM_DOUT_FILTERED[2]),
        .I4(I_MEM_DOUT_FILTERED[3]),
        .I5(I_MEM_DOUT_IBUF[31]),
        .O(\Q[98]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT5 #(
    .INIT(32'h20132033)) 
    \Q[98]_i_4 
       (.I0(I_MEM_DOUT_IBUF[2]),
        .I1(EX_BR_TAKEN),
        .I2(I_MEM_DOUT_IBUF[6]),
        .I3(I_MEM_DOUT_IBUF[4]),
        .I4(I_MEM_DOUT_IBUF[5]),
        .O(\Q[98]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[98]_i_5 
       (.I0(I_MEM_DOUT_IBUF[6]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[6]));
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \Q[98]_i_6 
       (.I0(I_MEM_DOUT_IBUF[3]),
        .I1(EX_BR_TAKEN),
        .O(I_MEM_DOUT_FILTERED[3]));
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \Q[99]_i_1 
       (.I0(\Q[109]_i_2_n_0 ),
        .I1(I_MEM_DOUT_IBUF[31]),
        .I2(CRF_RA2_OBUF[0]),
        .I3(\Q[123]_i_6_n_0 ),
        .O(ID_IMMEDIATE[20]));
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \Q[9]_i_1 
       (.I0(\custom_alu/fp32_add/significand_add0 [9]),
        .I1(\custom_alu/fp32_add/significand_add0 [24]),
        .I2(\custom_alu/fp32_add/significand_add0 [8]),
        .I3(\Q[30]_i_4__0_n_0 ),
        .O(\custom_alu/fp32_add/p_1_out [9]));
  LUT6 #(
    .INIT(64'h000007F7FFFF07F7)) 
    \Q[9]_i_10 
       (.I0(\Q[31]_i_13__0_n_0 ),
        .I1(\Q[29]_i_18__0_n_0 ),
        .I2(\Q[28]_i_20_n_0 ),
        .I3(\Q[17]_i_15_n_0 ),
        .I4(\Q[29]_i_10_n_0 ),
        .I5(\Q[35]_i_28_n_0 ),
        .O(\Q[9]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \Q[9]_i_10__0 
       (.I0(STALL_COUNTER_Q[5]),
        .I1(STALL_COUNTER_Q[4]),
        .I2(STALL_COUNTER_Q[3]),
        .O(\Q[9]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \Q[9]_i_11 
       (.I0(\Q[29]_i_7_n_0 ),
        .I1(EX_RF_RD1[27]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[153]),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(\custom_alu/int2fp/INT_VAL0 [27]),
        .O(\Q[9]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h9009090900000000)) 
    \Q[9]_i_11__0 
       (.I0(STALL_COUNTER_Q[1]),
        .I1(CUSTOM_INSTRUCTION_STALL_CYCLE[1]),
        .I2(STALL_COUNTER_Q[0]),
        .I3(\Q[112]_i_2_n_0 ),
        .I4(\Q[79]_i_3_n_0 ),
        .I5(\Q[9]_i_14_n_0 ),
        .O(\Q[9]_i_11__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF6FF6)) 
    \Q[9]_i_12 
       (.I0(CRF_RA2_OBUF[1]),
        .I1(ID_EX_Q[1]),
        .I2(CRF_RA2_OBUF[0]),
        .I3(ID_EX_Q[0]),
        .I4(\Q[9]_i_15_n_0 ),
        .O(\Q[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF01)) 
    \Q[9]_i_12__0 
       (.I0(\Q[31]_i_14__0_n_0 ),
        .I1(\Q[31]_i_10__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[67]_i_12_n_0 ),
        .I4(\Q[29]_i_7_n_0 ),
        .I5(\Q[35]_i_17_n_0 ),
        .O(\Q[9]_i_12__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF6FF6)) 
    \Q[9]_i_13 
       (.I0(CRF_RA1_OBUF[1]),
        .I1(ID_EX_Q[1]),
        .I2(CRF_RA1_OBUF[0]),
        .I3(ID_EX_Q[0]),
        .I4(\Q[9]_i_16_n_0 ),
        .O(\Q[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000DDDDDDD0DDD)) 
    \Q[9]_i_13__0 
       (.I0(ALU_DIN1[0]),
        .I1(\Q[21]_i_10__0_n_0 ),
        .I2(\Q[31]_i_11__0_n_0 ),
        .I3(\Q[47]_i_9_n_0 ),
        .I4(\Q[31]_i_14__0_n_0 ),
        .I5(\Q[35]_i_32_n_0 ),
        .O(\Q[9]_i_13__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT4 #(
    .INIT(16'h5559)) 
    \Q[9]_i_14 
       (.I0(STALL_COUNTER_Q[2]),
        .I1(\Q[31]_i_2_n_0 ),
        .I2(I_MEM_DOUT_IBUF[13]),
        .I3(I_MEM_DOUT_IBUF[14]),
        .O(\Q[9]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h6FF6)) 
    \Q[9]_i_15 
       (.I0(ID_EX_Q[2]),
        .I1(CRF_RA2_OBUF[2]),
        .I2(ID_EX_Q[3]),
        .I3(CRF_RA2_OBUF[3]),
        .O(\Q[9]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h6FF6)) 
    \Q[9]_i_16 
       (.I0(ID_EX_Q[2]),
        .I1(CRF_RA1_OBUF[2]),
        .I2(ID_EX_Q[3]),
        .I3(CRF_RA1_OBUF[3]),
        .O(\Q[9]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \Q[9]_i_1__0 
       (.I0(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[10] ),
        .I1(\Q[30]_i_2__1_n_0 ),
        .I2(\Q[9]_i_2_n_0 ),
        .I3(\Q[31]_i_2__1_n_0 ),
        .O(\custom_alu/FADD_Q [9]));
  LUT4 #(
    .INIT(16'hDDDF)) 
    \Q[9]_i_1__1 
       (.I0(RSTn_IBUF),
        .I1(LU_HAZARD),
        .I2(CUSTOM_EN),
        .I3(ID_WE_AFTER_LU3),
        .O(RST02_out));
  LUT6 #(
    .INIT(64'hFBAAFFFFFBAA0000)) 
    \Q[9]_i_1__2 
       (.I0(\Q[9]_i_2__0_n_0 ),
        .I1(\Q[9]_i_3__1_n_0 ),
        .I2(\Q[9]_i_4_n_0 ),
        .I3(\Q[34]_i_5_n_0 ),
        .I4(\FF_CUSTOM_EN/Q_reg_n_0_[0] ),
        .I5(D_MEM_ADDR_OBUF[4]),
        .O(data0[4]));
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \Q[9]_i_1__3 
       (.I0(\Q[9]_i_2__1_n_0 ),
        .I1(\Q[11]_i_3__0_n_0 ),
        .I2(\Q[9]_i_3__2_n_0 ),
        .I3(\Q[11]_i_5__1_n_0 ),
        .I4(MEM_D_MEM_ALU_FINAL1),
        .I5(EX_MEM_Q[9]),
        .O(data1[4]));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \Q[9]_i_2 
       (.I0(\custom_alu/fp32_add/sel0 [9]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .I2(\Q[9]_i_3__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [24]),
        .I4(\custom_alu/fp32_add/data23 [9]),
        .O(\Q[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[9]_i_2__0 
       (.I0(\custom_alu/MULT [4]),
        .I1(EX_CUSTOM_ALU_SEL[31]),
        .I2(\custom_alu/MULT [36]),
        .I3(EX_CUSTOM_ALU_SEL[30]),
        .I4(\custom_alu/Q [4]),
        .I5(EX_CUSTOM_ALU_SEL[29]),
        .O(\Q[9]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hF0AAFFCCF0AA00CC)) 
    \Q[9]_i_2__1 
       (.I0(D_MEM_DOUT_IBUF[12]),
        .I1(D_MEM_DOUT_IBUF[4]),
        .I2(D_MEM_DOUT_IBUF[28]),
        .I3(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I5(D_MEM_DOUT_IBUF[20]),
        .O(\Q[9]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00007FFF00008000)) 
    \Q[9]_i_2__2 
       (.I0(STALL_COUNTER_Q[8]),
        .I1(STALL_COUNTER_Q[6]),
        .I2(\Q[9]_i_4__1_n_0 ),
        .I3(STALL_COUNTER_Q[7]),
        .I4(STALL_COUNTER_D1),
        .I5(STALL_COUNTER_Q[9]),
        .O(STALL_COUNTER_D[9]));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'h40404000)) 
    \Q[9]_i_3 
       (.I0(D_MEM_CSN_OBUF),
        .I1(ID_EX_Q[124]),
        .I2(RSTn_IBUF),
        .I3(\stall_generator/LU_HAZARD1 ),
        .I4(\stall_generator/LU_HAZARD17_out ),
        .O(LU_HAZARD));
  LUT5 #(
    .INIT(32'hFF8B008B)) 
    \Q[9]_i_3__0 
       (.I0(\custom_alu/fp32_add/sel0 [7]),
        .I1(\custom_alu/fp32_add/sel0 [21]),
        .I2(\Q[9]_i_4__0_n_0 ),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(\custom_alu/fp32_add/sel0 [8]),
        .O(\Q[9]_i_3__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \Q[9]_i_3__1 
       (.I0(\Q[65]_i_5_n_0 ),
        .I1(\custom_alu/fp32_mult/product_mantissa [4]),
        .O(\Q[9]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \Q[9]_i_3__2 
       (.I0(D_MEM_DOUT_IBUF[4]),
        .I1(D_MEM_DOUT_IBUF[20]),
        .I2(\FF_EX_MEM_TEMP/Q_reg_n_0_[0] ),
        .I3(D_MEM_DOUT_IBUF[28]),
        .I4(\FF_EX_MEM_TEMP/Q_reg_n_0_[1] ),
        .I5(D_MEM_DOUT_IBUF[12]),
        .O(\Q[9]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h2222202220202020)) 
    \Q[9]_i_4 
       (.I0(\Q[9]_i_5__0_n_0 ),
        .I1(\Q[9]_i_6__1_n_0 ),
        .I2(EX_CUSTOM_ALU_SEL[27]),
        .I3(\Q[9]_i_7__0_n_0 ),
        .I4(\Q[9]_i_8__0_n_0 ),
        .I5(EX_CUSTOM_ALU_SEL[26]),
        .O(\Q[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[9]_i_4__0 
       (.I0(\custom_alu/fp32_add/sel0 [6]),
        .I1(\custom_alu/fp32_add/sel0 [20]),
        .I2(\custom_alu/fp32_add/sel0 [5]),
        .I3(\custom_alu/fp32_add/sel0 [19]),
        .I4(\Q[9]_i_5_n_0 ),
        .O(\Q[9]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \Q[9]_i_4__1 
       (.I0(STALL_COUNTER_Q[5]),
        .I1(STALL_COUNTER_Q[3]),
        .I2(STALL_COUNTER_Q[1]),
        .I3(STALL_COUNTER_Q[0]),
        .I4(STALL_COUNTER_Q[2]),
        .I5(STALL_COUNTER_Q[4]),
        .O(\Q[9]_i_4__1_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \Q[9]_i_5 
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [17]),
        .I4(\Q[9]_i_6__0_n_0 ),
        .O(\Q[9]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0047FFFFFFFF)) 
    \Q[9]_i_5__0 
       (.I0(INT0_carry_i_10_n_0),
        .I1(ALU_DIN1[23]),
        .I2(INT0_carry_i_9_n_0),
        .I3(INT0_carry_i_6_n_0),
        .I4(PSUM3__0_carry__0_i_10__2_n_0),
        .I5(EX_CUSTOM_ALU_SEL[27]),
        .O(\Q[9]_i_5__0_n_0 ));
  LUT5 #(
    .INIT(32'h00009009)) 
    \Q[9]_i_6 
       (.I0(CUSTOM_RS2),
        .I1(EX_CUSTOM_RD),
        .I2(CRF_RA2_OBUF[4]),
        .I3(ID_EX_Q[4]),
        .I4(\Q[9]_i_12_n_0 ),
        .O(\stall_generator/LU_HAZARD1 ));
  LUT6 #(
    .INIT(64'h4744477747774777)) 
    \Q[9]_i_6__0 
       (.I0(\custom_alu/fp32_add/sel0 [2]),
        .I1(\custom_alu/fp32_add/sel0 [16]),
        .I2(\custom_alu/fp32_add/sel0 [1]),
        .I3(\custom_alu/fp32_add/sel0 [15]),
        .I4(\custom_alu/fp32_add/sel0 [0]),
        .I5(\custom_alu/fp32_add/sel0 [14]),
        .O(\Q[9]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAEAAAA)) 
    \Q[9]_i_6__1 
       (.I0(EX_CUSTOM_ALU_SEL[28]),
        .I1(EX_RF_RD1[31]),
        .I2(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I3(ID_EX_Q[157]),
        .I4(EX_CUSTOM_ALU_SEL[27]),
        .I5(\custom_alu/fp2int/INT0 [4]),
        .O(\Q[9]_i_6__1_n_0 ));
  LUT5 #(
    .INIT(32'h00009009)) 
    \Q[9]_i_7 
       (.I0(CUSTOM_RS1),
        .I1(EX_CUSTOM_RD),
        .I2(CRF_RA1_OBUF[4]),
        .I3(ID_EX_Q[4]),
        .I4(\Q[9]_i_13_n_0 ),
        .O(\stall_generator/LU_HAZARD17_out ));
  LUT6 #(
    .INIT(64'h54545400FFFFFFFF)) 
    \Q[9]_i_7__0 
       (.I0(\Q[9]_i_9_n_0 ),
        .I1(\Q[9]_i_10_n_0 ),
        .I2(\Q[9]_i_11_n_0 ),
        .I3(\Q[9]_i_12__0_n_0 ),
        .I4(\Q[9]_i_13__0_n_0 ),
        .I5(\Q[26]_i_7_n_0 ),
        .O(\Q[9]_i_7__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \Q[9]_i_8 
       (.I0(STALL_COUNTER_Q[9]),
        .O(\Q[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \Q[9]_i_8__0 
       (.I0(\Q[35]_i_19_n_0 ),
        .I1(\Q[28]_i_6_n_0 ),
        .I2(\Q[35]_i_21_n_0 ),
        .I3(\Q[35]_i_18_n_0 ),
        .I4(\Q[35]_i_22_n_0 ),
        .I5(\Q[35]_i_16_n_0 ),
        .O(\Q[9]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hBB8BB888B888B888)) 
    \Q[9]_i_9 
       (.I0(\Q[35]_i_27_n_0 ),
        .I1(\Q[35]_i_17_n_0 ),
        .I2(\Q[28]_i_12_n_0 ),
        .I3(\Q[35]_i_26_n_0 ),
        .I4(\Q[35]_i_29_n_0 ),
        .I5(\Q[23]_i_13__0_n_0 ),
        .O(\Q[9]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \Q[9]_i_9__0 
       (.I0(STALL_COUNTER_Q[8]),
        .I1(STALL_COUNTER_Q[7]),
        .I2(STALL_COUNTER_Q[6]),
        .O(\Q[9]_i_9__0_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[12]_i_1 
       (.CI(\Q_reg[8]_i_1_n_0 ),
        .CO({\Q_reg[12]_i_1_n_0 ,\Q_reg[12]_i_1_n_1 ,\Q_reg[12]_i_1_n_2 ,\Q_reg[12]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(IF_PC_ADD4[12:9]),
        .S({\Q[12]_i_2__1_n_0 ,\Q[12]_i_3__3_n_0 ,\Q[12]_i_4__2_n_0 ,\Q[12]_i_5__1_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[12]_i_10 
       (.CI(\Q_reg[49]_i_6_n_0 ),
        .CO({\Q_reg[12]_i_10_n_0 ,\Q_reg[12]_i_10_n_1 ,\Q_reg[12]_i_10_n_2 ,\Q_reg[12]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_mult/product_mantissa [7:4]),
        .S({\Q[12]_i_14_n_0 ,\Q[12]_i_15__0_n_0 ,\Q[12]_i_16__0_n_0 ,\Q[12]_i_17__0_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[12]_i_2 
       (.CI(\Q_reg[8]_i_2_n_0 ),
        .CO({\Q_reg[12]_i_2_n_0 ,\Q_reg[12]_i_2_n_1 ,\Q_reg[12]_i_2_n_2 ,\Q_reg[12]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/data23 [12:9]),
        .S({\Q[12]_i_4__0_n_0 ,\Q[12]_i_5__0_n_0 ,\Q[12]_i_6__0_n_0 ,\Q[12]_i_7_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[12]_i_2__0 
       (.CI(\Q_reg[8]_i_2__0_n_0 ),
        .CO({\Q_reg[12]_i_2__0_n_0 ,\Q_reg[12]_i_2__0_n_1 ,\Q_reg[12]_i_2__0_n_2 ,\Q_reg[12]_i_2__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_b_add_sub [11:8]),
        .O(\custom_alu/fp32_add/significand_add0 [11:8]),
        .S({\fp32_add/Q[12]_i_7_n_0 ,\fp32_add/Q[12]_i_8_n_0 ,\fp32_add/Q[12]_i_9_n_0 ,\fp32_add/Q[12]_i_10_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[16]_i_1 
       (.CI(\Q_reg[12]_i_1_n_0 ),
        .CO({\Q_reg[16]_i_1_n_0 ,\Q_reg[16]_i_1_n_1 ,\Q_reg[16]_i_1_n_2 ,\Q_reg[16]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(IF_PC_ADD4[16:13]),
        .S({\Q[16]_i_2__3_n_0 ,\Q[16]_i_3__3_n_0 ,\Q[16]_i_4__2_n_0 ,\Q[16]_i_5__1_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[16]_i_13 
       (.CI(\Q_reg[49]_i_18_n_0 ),
        .CO({\Q_reg[16]_i_13_n_0 ,\Q_reg[16]_i_13_n_1 ,\Q_reg[16]_i_13_n_2 ,\Q_reg[16]_i_13_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/p_1_in [34:31]),
        .O({\Q_reg[16]_i_13_n_4 ,\Q_reg[16]_i_13_n_5 ,\Q_reg[16]_i_13_n_6 ,\Q_reg[16]_i_13_n_7 }),
        .S({\fp32_mult/mult24_0/Q[16]_i_14_n_0 ,\fp32_mult/mult24_0/Q[16]_i_15_n_0 ,\fp32_mult/mult24_0/Q[16]_i_16_n_0 ,\fp32_mult/mult24_0/Q[16]_i_17_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[16]_i_2 
       (.CI(\Q_reg[12]_i_2__0_n_0 ),
        .CO({\Q_reg[16]_i_2_n_0 ,\Q_reg[16]_i_2_n_1 ,\Q_reg[16]_i_2_n_2 ,\Q_reg[16]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_b_add_sub [15:12]),
        .O(\custom_alu/fp32_add/significand_add0 [15:12]),
        .S({\fp32_add/Q[16]_i_7_n_0 ,\fp32_add/Q[16]_i_8_n_0 ,\fp32_add/Q[16]_i_9_n_0 ,\fp32_add/Q[16]_i_10_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[16]_i_5 
       (.CI(\Q_reg[12]_i_2_n_0 ),
        .CO({\Q_reg[16]_i_5_n_0 ,\Q_reg[16]_i_5_n_1 ,\Q_reg[16]_i_5_n_2 ,\Q_reg[16]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/data23 [16:13]),
        .S({\Q[16]_i_7_n_0 ,\Q[16]_i_8_n_0 ,\Q[16]_i_9_n_0 ,\Q[16]_i_10_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[16]_i_6 
       (.CI(\Q_reg[12]_i_10_n_0 ),
        .CO({\Q_reg[16]_i_6_n_0 ,\Q_reg[16]_i_6_n_1 ,\Q_reg[16]_i_6_n_2 ,\Q_reg[16]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_mult/product_mantissa [11:8]),
        .S({\Q[16]_i_9__0_n_0 ,\Q[16]_i_10__0_n_0 ,\Q[16]_i_11__1_n_0 ,\Q[16]_i_12__1_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_10 
       (.CI(\Q_reg[171]_i_16_n_0 ),
        .CO({\branch_comp/LT20_in ,\Q_reg[171]_i_10_n_1 ,\Q_reg[171]_i_10_n_2 ,\Q_reg[171]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_17_n_0 ,\Q[171]_i_18_n_0 ,\Q[171]_i_19_n_0 ,\Q[171]_i_20_n_0 }),
        .S({\Q[171]_i_21_n_0 ,\Q[171]_i_22_n_0 ,\Q[171]_i_23_n_0 ,\Q[171]_i_24_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_11 
       (.CI(\Q_reg[171]_i_25_n_0 ),
        .CO({\Q_reg[171]_i_11_n_0 ,\Q_reg[171]_i_11_n_1 ,\Q_reg[171]_i_11_n_2 ,\Q_reg[171]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_26_n_0 ,\Q[171]_i_27_n_0 ,\Q[171]_i_28_n_0 ,\Q[171]_i_29_n_0 }),
        .S({\Q[171]_i_30_n_0 ,\Q[171]_i_31_n_0 ,\Q[171]_i_32_n_0 ,\Q[171]_i_33_n_0 }));
  CARRY4 \Q_reg[171]_i_12 
       (.CI(\Q_reg[171]_i_34_n_0 ),
        .CO({\Q_reg[171]_i_12_n_0 ,\Q_reg[171]_i_12_n_1 ,\Q_reg[171]_i_12_n_2 ,\Q_reg[171]_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\Q[171]_i_35_n_0 ,\Q[171]_i_36_n_0 ,\Q[171]_i_37_n_0 ,\Q[171]_i_38_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_16 
       (.CI(\Q_reg[171]_i_39_n_0 ),
        .CO({\Q_reg[171]_i_16_n_0 ,\Q_reg[171]_i_16_n_1 ,\Q_reg[171]_i_16_n_2 ,\Q_reg[171]_i_16_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_40_n_0 ,\Q[171]_i_41_n_0 ,\Q[171]_i_42_n_0 ,\Q[171]_i_43_n_0 }),
        .S({\Q[171]_i_44_n_0 ,\Q[171]_i_45_n_0 ,\Q[171]_i_46_n_0 ,\Q[171]_i_47_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_25 
       (.CI(\Q_reg[171]_i_48_n_0 ),
        .CO({\Q_reg[171]_i_25_n_0 ,\Q_reg[171]_i_25_n_1 ,\Q_reg[171]_i_25_n_2 ,\Q_reg[171]_i_25_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_49_n_0 ,\Q[171]_i_50_n_0 ,\Q[171]_i_51_n_0 ,\Q[171]_i_52_n_0 }),
        .S({\Q[171]_i_53_n_0 ,\Q[171]_i_54_n_0 ,\Q[171]_i_55_n_0 ,\Q[171]_i_56_n_0 }));
  CARRY4 \Q_reg[171]_i_34 
       (.CI(\<const0> ),
        .CO({\Q_reg[171]_i_34_n_0 ,\Q_reg[171]_i_34_n_1 ,\Q_reg[171]_i_34_n_2 ,\Q_reg[171]_i_34_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\Q[171]_i_57_n_0 ,\Q[171]_i_58_n_0 ,\Q[171]_i_59_n_0 ,\Q[171]_i_60_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_39 
       (.CI(\Q_reg[171]_i_63_n_0 ),
        .CO({\Q_reg[171]_i_39_n_0 ,\Q_reg[171]_i_39_n_1 ,\Q_reg[171]_i_39_n_2 ,\Q_reg[171]_i_39_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_64_n_0 ,\Q[171]_i_65_n_0 ,\Q[171]_i_66_n_0 ,\Q[171]_i_67_n_0 }),
        .S({\Q[171]_i_68_n_0 ,\Q[171]_i_69_n_0 ,\Q[171]_i_70_n_0 ,\Q[171]_i_71_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_48 
       (.CI(\Q_reg[171]_i_73_n_0 ),
        .CO({\Q_reg[171]_i_48_n_0 ,\Q_reg[171]_i_48_n_1 ,\Q_reg[171]_i_48_n_2 ,\Q_reg[171]_i_48_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_64_n_0 ,\Q[171]_i_74_n_0 ,\Q[171]_i_75_n_0 ,\Q[171]_i_76_n_0 }),
        .S({\Q[171]_i_77_n_0 ,\Q[171]_i_78_n_0 ,\Q[171]_i_79_n_0 ,\Q[171]_i_80_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_63 
       (.CI(\<const0> ),
        .CO({\Q_reg[171]_i_63_n_0 ,\Q_reg[171]_i_63_n_1 ,\Q_reg[171]_i_63_n_2 ,\Q_reg[171]_i_63_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_85_n_0 ,\Q[171]_i_86_n_0 ,\Q[171]_i_87_n_0 ,\Q[171]_i_88_n_0 }),
        .S({\Q[171]_i_89_n_0 ,\Q[171]_i_90_n_0 ,\Q[171]_i_91_n_0 ,\Q[171]_i_92_n_0 }));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \Q_reg[171]_i_73 
       (.CI(\<const0> ),
        .CO({\Q_reg[171]_i_73_n_0 ,\Q_reg[171]_i_73_n_1 ,\Q_reg[171]_i_73_n_2 ,\Q_reg[171]_i_73_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\Q[171]_i_93_n_0 ,\Q[171]_i_94_n_0 ,\Q[171]_i_95_n_0 ,\Q[171]_i_96_n_0 }),
        .S({\Q[171]_i_97_n_0 ,\Q[171]_i_98_n_0 ,\Q[171]_i_99_n_0 ,\Q[171]_i_100_n_0 }));
  CARRY4 \Q_reg[171]_i_8 
       (.CI(\Q_reg[171]_i_12_n_0 ),
        .CO({\branch_comp/EQ ,\Q_reg[171]_i_8_n_2 ,\Q_reg[171]_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\Q[171]_i_13_n_0 ,\Q[171]_i_14_n_0 ,\Q[171]_i_15_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[20]_i_1 
       (.CI(\Q_reg[16]_i_1_n_0 ),
        .CO({\Q_reg[20]_i_1_n_0 ,\Q_reg[20]_i_1_n_1 ,\Q_reg[20]_i_1_n_2 ,\Q_reg[20]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(IF_PC_ADD4[20:17]),
        .S({\Q[20]_i_2__3_n_0 ,\Q[20]_i_3__4_n_0 ,\Q[20]_i_4__3_n_0 ,\Q[20]_i_5__2_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[20]_i_2 
       (.CI(\Q_reg[16]_i_2_n_0 ),
        .CO({\Q_reg[20]_i_2_n_0 ,\Q_reg[20]_i_2_n_1 ,\Q_reg[20]_i_2_n_2 ,\Q_reg[20]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_b_add_sub [19:16]),
        .O(\custom_alu/fp32_add/significand_add0 [19:16]),
        .S({\fp32_add/Q[20]_i_7_n_0 ,\fp32_add/Q[20]_i_8_n_0 ,\fp32_add/Q[20]_i_9_n_0 ,\fp32_add/Q[20]_i_10_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[20]_i_6 
       (.CI(\Q_reg[16]_i_6_n_0 ),
        .CO({\Q_reg[20]_i_6_n_0 ,\Q_reg[20]_i_6_n_1 ,\Q_reg[20]_i_6_n_2 ,\Q_reg[20]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_mult/product_mantissa [15:12]),
        .S({\Q[20]_i_9__0_n_0 ,\Q[20]_i_10__0_n_0 ,\Q[20]_i_11__0_n_0 ,\Q[20]_i_12__0_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[22]_i_2 
       (.CI(\Q_reg[22]_i_4_n_0 ),
        .CO(\Q_reg[22]_i_2_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/data23 [22:21]),
        .S({\<const0> ,\<const0> ,\Q[22]_i_5_n_0 ,\Q[22]_i_6_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[22]_i_4 
       (.CI(\Q_reg[16]_i_5_n_0 ),
        .CO({\Q_reg[22]_i_4_n_0 ,\Q_reg[22]_i_4_n_1 ,\Q_reg[22]_i_4_n_2 ,\Q_reg[22]_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/data23 [20:17]),
        .S({\Q[22]_i_8_n_0 ,\Q[22]_i_9_n_0 ,\Q[22]_i_10_n_0 ,\Q[22]_i_11_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[23]_i_2 
       (.CI(\Q_reg[20]_i_2_n_0 ),
        .CO({\Q_reg[23]_i_2_n_0 ,\Q_reg[23]_i_2_n_1 ,\Q_reg[23]_i_2_n_2 ,\Q_reg[23]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_b_add_sub [23:20]),
        .O(\custom_alu/fp32_add/significand_add0 [23:20]),
        .S({\Q[23]_i_7__0_n_0 ,\fp32_add/Q[23]_i_8_n_0 ,\fp32_add/Q[23]_i_9_n_0 ,\fp32_add/Q[23]_i_10_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[24]_i_1 
       (.CI(\Q_reg[20]_i_1_n_0 ),
        .CO({\Q_reg[24]_i_1_n_0 ,\Q_reg[24]_i_1_n_1 ,\Q_reg[24]_i_1_n_2 ,\Q_reg[24]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(IF_PC_ADD4[24:21]),
        .S({\Q[24]_i_2__1_n_0 ,\Q[24]_i_3__0_n_0 ,\Q[24]_i_4__1_n_0 ,\Q[24]_i_5__0_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[27]_i_8 
       (.CI(\Q_reg[65]_i_6_n_0 ),
        .CO({\Q_reg[27]_i_8_n_2 ,\Q_reg[27]_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_mult/product_mantissa [22:20]),
        .S({\<const0> ,\Q[27]_i_16_n_0 ,\Q[27]_i_17_n_0 ,\Q[27]_i_18_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[28]_i_1 
       (.CI(\Q_reg[24]_i_1_n_0 ),
        .CO({\Q_reg[28]_i_1_n_0 ,\Q_reg[28]_i_1_n_1 ,\Q_reg[28]_i_1_n_2 ,\Q_reg[28]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(IF_PC_ADD4[28:25]),
        .S({\Q[28]_i_2__1_n_0 ,\Q[28]_i_3__0_n_0 ,\Q[28]_i_4__0_n_0 ,\Q[28]_i_5__0_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[29]_i_14 
       (.CI(\Q_reg[29]_i_9_n_0 ),
        .CO({\Q_reg[29]_i_14_n_0 ,\Q_reg[29]_i_14_n_1 ,\Q_reg[29]_i_14_n_2 ,\Q_reg[29]_i_14_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [28:25]),
        .S({\Q[29]_i_23_n_0 ,\Q[29]_i_24_n_0 ,\Q[29]_i_25_n_0 ,\Q[29]_i_26_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[29]_i_9 
       (.CI(\Q_reg[30]_i_18_n_0 ),
        .CO({\Q_reg[29]_i_9_n_0 ,\Q_reg[29]_i_9_n_1 ,\Q_reg[29]_i_9_n_2 ,\Q_reg[29]_i_9_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [24:21]),
        .S({\Q[29]_i_15_n_0 ,\Q[29]_i_16_n_0 ,\custom_alu/int2fp/INT_VAL1 [22:21]}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[30]_i_18 
       (.CI(\Q_reg[35]_i_31_n_0 ),
        .CO({\Q_reg[30]_i_18_n_0 ,\Q_reg[30]_i_18_n_1 ,\Q_reg[30]_i_18_n_2 ,\Q_reg[30]_i_18_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [20:17]),
        .S({\custom_alu/int2fp/INT_VAL1 [20:18],\Q[30]_i_22_n_0 }));
  CARRY4 \Q_reg[30]_i_3 
       (.CI(\Q_reg[23]_i_2_n_0 ),
        .CO(\custom_alu/fp32_add/significand_add0 [24]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[30]_i_7 
       (.CI(\Q_reg[29]_i_14_n_0 ),
        .CO(\Q_reg[30]_i_7_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [30:29]),
        .S({\<const0> ,\<const0> ,\Q[30]_i_11_n_0 ,\Q[30]_i_12_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[31]_i_1 
       (.CI(\Q_reg[28]_i_1_n_0 ),
        .CO({\Q_reg[31]_i_1_n_2 ,\Q_reg[31]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(IF_PC_ADD4[31:29]),
        .S({\<const0> ,\Q[31]_i_2__4_n_0 ,\Q[31]_i_3__3_n_0 ,\Q[31]_i_4__2_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[35]_i_30 
       (.CI(\Q_reg[35]_i_34_n_0 ),
        .CO({\Q_reg[35]_i_30_n_0 ,\Q_reg[35]_i_30_n_1 ,\Q_reg[35]_i_30_n_2 ,\Q_reg[35]_i_30_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [12:9]),
        .S({\Q[35]_i_35_n_0 ,\Q[35]_i_36_n_0 ,\Q[35]_i_37_n_0 ,\Q[35]_i_38_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[35]_i_31 
       (.CI(\Q_reg[35]_i_30_n_0 ),
        .CO({\Q_reg[35]_i_31_n_0 ,\Q_reg[35]_i_31_n_1 ,\Q_reg[35]_i_31_n_2 ,\Q_reg[35]_i_31_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [16:13]),
        .S({\Q[35]_i_39_n_0 ,\Q[35]_i_40_n_0 ,\Q[35]_i_41_n_0 ,\Q[35]_i_42_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[35]_i_33 
       (.CI(\<const0> ),
        .CO({\Q_reg[35]_i_33_n_0 ,\Q_reg[35]_i_33_n_1 ,\Q_reg[35]_i_33_n_2 ,\Q_reg[35]_i_33_n_3 }),
        .CYINIT(\custom_alu/int2fp/INT_VAL1 [0]),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [4:1]),
        .S(\custom_alu/int2fp/INT_VAL1 [4:1]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[35]_i_34 
       (.CI(\Q_reg[35]_i_33_n_0 ),
        .CO({\Q_reg[35]_i_34_n_0 ,\Q_reg[35]_i_34_n_1 ,\Q_reg[35]_i_34_n_2 ,\Q_reg[35]_i_34_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/int2fp/INT_VAL0 [8:5]),
        .S({\Q[35]_i_48_n_0 ,\custom_alu/int2fp/INT_VAL1 [7:5]}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[49]_i_17 
       (.CI(\Q_reg[49]_i_21_n_0 ),
        .CO({\Q_reg[49]_i_17_n_0 ,\Q_reg[49]_i_17_n_1 ,\Q_reg[49]_i_17_n_2 ,\Q_reg[49]_i_17_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/p_1_in [26:23]),
        .O({\Q_reg[49]_i_17_n_4 ,\Q_reg[49]_i_17_n_5 ,\Q_reg[49]_i_17_n_6 ,\Q_reg[49]_i_17_n_7 }),
        .S({\fp32_mult/mult24_0/Q[49]_i_24_n_0 ,\fp32_mult/mult24_0/Q[49]_i_25_n_0 ,\fp32_mult/mult24_0/Q[49]_i_26_n_0 ,\fp32_mult/mult24_0/Q[49]_i_27_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[49]_i_18 
       (.CI(\Q_reg[49]_i_17_n_0 ),
        .CO({\Q_reg[49]_i_18_n_0 ,\Q_reg[49]_i_18_n_1 ,\Q_reg[49]_i_18_n_2 ,\Q_reg[49]_i_18_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/p_1_in [30:27]),
        .O({\Q_reg[49]_i_18_n_4 ,\Q_reg[49]_i_18_n_5 ,\Q_reg[49]_i_18_n_6 ,\Q_reg[49]_i_18_n_7 }),
        .S({\fp32_mult/mult24_0/Q[49]_i_28_n_0 ,\fp32_mult/mult24_0/Q[49]_i_29_n_0 ,\fp32_mult/mult24_0/Q[49]_i_30_n_0 ,\fp32_mult/mult24_0/Q[49]_i_31_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[49]_i_21 
       (.CI(\Q_reg[49]_i_35_n_0 ),
        .CO({\Q_reg[49]_i_21_n_0 ,\Q_reg[49]_i_21_n_1 ,\Q_reg[49]_i_21_n_2 ,\Q_reg[49]_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/p_1_in [22:19]),
        .O({\Q_reg[49]_i_21_n_4 ,\Q_reg[49]_i_21_n_5 ,\Q_reg[49]_i_21_n_6 ,\Q_reg[49]_i_21_n_7 }),
        .S({\fp32_mult/mult24_0/Q[49]_i_37_n_0 ,\fp32_mult/mult24_0/Q[49]_i_38_n_0 ,\fp32_mult/mult24_0/Q[49]_i_39_n_0 ,\fp32_mult/mult24_0/Q[49]_i_40_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[49]_i_32 
       (.CI(\<const0> ),
        .CO({\Q_reg[49]_i_32_n_0 ,\Q_reg[49]_i_32_n_1 ,\Q_reg[49]_i_32_n_2 ,\Q_reg[49]_i_32_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/fp32_mult/p_1_in [14:12],\<const0> }),
        .O({\Q_reg[49]_i_32_n_4 ,\Q_reg[49]_i_32_n_5 ,\Q_reg[49]_i_32_n_6 ,\Q_reg[49]_i_32_n_7 }),
        .S({\fp32_mult/mult24_0/Q[49]_i_41_n_0 ,\fp32_mult/mult24_0/Q[49]_i_42_n_0 ,\fp32_mult/mult24_0/Q[49]_i_43_n_0 ,\custom_alu/fp32_mult/p_1_in [11]}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[49]_i_35 
       (.CI(\Q_reg[49]_i_32_n_0 ),
        .CO({\Q_reg[49]_i_35_n_0 ,\Q_reg[49]_i_35_n_1 ,\Q_reg[49]_i_35_n_2 ,\Q_reg[49]_i_35_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/p_1_in [18:15]),
        .O({\Q_reg[49]_i_35_n_4 ,\Q_reg[49]_i_35_n_5 ,\Q_reg[49]_i_35_n_6 ,\Q_reg[49]_i_35_n_7 }),
        .S({\fp32_mult/mult24_0/Q[49]_i_44_n_0 ,\fp32_mult/mult24_0/Q[49]_i_45_n_0 ,\fp32_mult/mult24_0/Q[49]_i_46_n_0 ,\fp32_mult/mult24_0/Q[49]_i_47_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[49]_i_6 
       (.CI(\<const0> ),
        .CO({\Q_reg[49]_i_6_n_0 ,\Q_reg[49]_i_6_n_1 ,\Q_reg[49]_i_6_n_2 ,\Q_reg[49]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\Q[49]_i_11_n_0 }),
        .O(\custom_alu/fp32_mult/product_mantissa [3:0]),
        .S({\Q[49]_i_12_n_0 ,\Q[49]_i_13_n_0 ,\Q[49]_i_14_n_0 ,\Q[49]_i_15_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[4]_i_1 
       (.CI(\<const0> ),
        .CO({\Q_reg[4]_i_1_n_0 ,\Q_reg[4]_i_1_n_1 ,\Q_reg[4]_i_1_n_2 ,\Q_reg[4]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const1> ,\<const0> }),
        .O(IF_PC_ADD4[4:1]),
        .S({\Q[4]_i_2_n_0 ,\Q[4]_i_3__1_n_0 ,\Q[4]_i_4__1_n_0 ,\Q[4]_i_5__1_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[4]_i_2 
       (.CI(\<const0> ),
        .CO({\Q_reg[4]_i_2_n_0 ,\Q_reg[4]_i_2_n_1 ,\Q_reg[4]_i_2_n_2 ,\Q_reg[4]_i_2_n_3 }),
        .CYINIT(\Q[4]_i_4__0_n_0 ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/data23 [4:1]),
        .S({\Q[4]_i_5__0_n_0 ,\Q[4]_i_6__0_n_0 ,\Q[4]_i_7_n_0 ,\Q[4]_i_8_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[4]_i_2__0 
       (.CI(\<const0> ),
        .CO({\Q_reg[4]_i_2__0_n_0 ,\Q_reg[4]_i_2__0_n_1 ,\Q_reg[4]_i_2__0_n_2 ,\Q_reg[4]_i_2__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_b_add_sub [3:0]),
        .O(\custom_alu/fp32_add/significand_add0 [3:0]),
        .S({\fp32_add/Q[4]_i_7_n_0 ,\fp32_add/Q[4]_i_8_n_0 ,\fp32_add/Q[4]_i_9_n_0 ,\fp32_add/Q[4]_i_10_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[65]_i_6 
       (.CI(\Q_reg[20]_i_6_n_0 ),
        .CO({\Q_reg[65]_i_6_n_0 ,\Q_reg[65]_i_6_n_1 ,\Q_reg[65]_i_6_n_2 ,\Q_reg[65]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_mult/product_mantissa [19:16]),
        .S({\Q[65]_i_9_n_0 ,\Q[65]_i_10_n_0 ,\Q[65]_i_11_n_0 ,\Q[65]_i_12_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[67]_i_2 
       (.CI(\<const0> ),
        .CO({\Q_reg[67]_i_2_n_0 ,\Q_reg[67]_i_2_n_1 ,\Q_reg[67]_i_2_n_2 ,\Q_reg[67]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_sub_complement [3:0]),
        .O(\custom_alu/fp32_add/significand_sub0 [3:0]),
        .S({\fp32_add/Q[67]_i_4_n_0 ,\fp32_add/Q[67]_i_5_n_0 ,\fp32_add/Q[67]_i_6_n_0 ,\fp32_add/Q[67]_i_7_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[67]_i_3 
       (.CI(\<const0> ),
        .CO({\Q_reg[67]_i_3_n_0 ,\Q_reg[67]_i_3_n_1 ,\Q_reg[67]_i_3_n_2 ,\Q_reg[67]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\custom_alu/fp32_add/significand_sub_complement1 }),
        .O(\custom_alu/fp32_add/significand_sub_complement [3:0]),
        .S({\Q[67]_i_9_n_0 ,\Q[67]_i_10_n_0 ,\Q[67]_i_11_n_0 ,\Q[67]_i_12__0_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[71]_i_2 
       (.CI(\Q_reg[67]_i_2_n_0 ),
        .CO({\Q_reg[71]_i_2_n_0 ,\Q_reg[71]_i_2_n_1 ,\Q_reg[71]_i_2_n_2 ,\Q_reg[71]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_sub_complement [7:4]),
        .O(\custom_alu/fp32_add/significand_sub0 [7:4]),
        .S({\fp32_add/Q[71]_i_4_n_0 ,\fp32_add/Q[71]_i_5_n_0 ,\fp32_add/Q[71]_i_6_n_0 ,\fp32_add/Q[71]_i_7_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[71]_i_3 
       (.CI(\Q_reg[67]_i_3_n_0 ),
        .CO({\Q_reg[71]_i_3_n_0 ,\Q_reg[71]_i_3_n_1 ,\Q_reg[71]_i_3_n_2 ,\Q_reg[71]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/significand_sub_complement [7:4]),
        .S({\Q[71]_i_8_n_0 ,\Q[71]_i_9_n_0 ,\Q[71]_i_10_n_0 ,\Q[71]_i_11_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[75]_i_2 
       (.CI(\Q_reg[71]_i_2_n_0 ),
        .CO({\Q_reg[75]_i_2_n_0 ,\Q_reg[75]_i_2_n_1 ,\Q_reg[75]_i_2_n_2 ,\Q_reg[75]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_sub_complement [11:8]),
        .O(\custom_alu/fp32_add/significand_sub0 [11:8]),
        .S({\fp32_add/Q[75]_i_4_n_0 ,\fp32_add/Q[75]_i_5_n_0 ,\fp32_add/Q[75]_i_6_n_0 ,\fp32_add/Q[75]_i_7_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[75]_i_3 
       (.CI(\Q_reg[71]_i_3_n_0 ),
        .CO({\Q_reg[75]_i_3_n_0 ,\Q_reg[75]_i_3_n_1 ,\Q_reg[75]_i_3_n_2 ,\Q_reg[75]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/significand_sub_complement [11:8]),
        .S({\Q[75]_i_8_n_0 ,\Q[75]_i_9_n_0 ,\Q[75]_i_10_n_0 ,\Q[75]_i_11_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[79]_i_2 
       (.CI(\Q_reg[75]_i_2_n_0 ),
        .CO({\Q_reg[79]_i_2_n_0 ,\Q_reg[79]_i_2_n_1 ,\Q_reg[79]_i_2_n_2 ,\Q_reg[79]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_sub_complement [15:12]),
        .O(\custom_alu/fp32_add/significand_sub0 [15:12]),
        .S({\fp32_add/Q[79]_i_4_n_0 ,\fp32_add/Q[79]_i_5_n_0 ,\fp32_add/Q[79]_i_6_n_0 ,\fp32_add/Q[79]_i_7_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[79]_i_3 
       (.CI(\Q_reg[75]_i_3_n_0 ),
        .CO({\Q_reg[79]_i_3_n_0 ,\Q_reg[79]_i_3_n_1 ,\Q_reg[79]_i_3_n_2 ,\Q_reg[79]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/significand_sub_complement [15:12]),
        .S({\Q[79]_i_8_n_0 ,\Q[79]_i_9_n_0 ,\Q[79]_i_10_n_0 ,\Q[79]_i_11_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[83]_i_2 
       (.CI(\Q_reg[79]_i_2_n_0 ),
        .CO({\Q_reg[83]_i_2_n_0 ,\Q_reg[83]_i_2_n_1 ,\Q_reg[83]_i_2_n_2 ,\Q_reg[83]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_sub_complement [19:16]),
        .O(\custom_alu/fp32_add/significand_sub0 [19:16]),
        .S({\fp32_add/Q[83]_i_4_n_0 ,\fp32_add/Q[83]_i_5_n_0 ,\fp32_add/Q[83]_i_6_n_0 ,\fp32_add/Q[83]_i_7_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[83]_i_3 
       (.CI(\Q_reg[79]_i_3_n_0 ),
        .CO({\Q_reg[83]_i_3_n_0 ,\Q_reg[83]_i_3_n_1 ,\Q_reg[83]_i_3_n_2 ,\Q_reg[83]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/significand_sub_complement [19:16]),
        .S({\Q[83]_i_8_n_0 ,\Q[83]_i_9_n_0 ,\Q[83]_i_10_n_0 ,\Q[83]_i_11_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[87]_i_2 
       (.CI(\Q_reg[83]_i_2_n_0 ),
        .CO({\Q_reg[87]_i_2_n_0 ,\Q_reg[87]_i_2_n_1 ,\Q_reg[87]_i_2_n_2 ,\Q_reg[87]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_sub_complement [23:20]),
        .O(\custom_alu/fp32_add/significand_sub0 [23:20]),
        .S({\Q[87]_i_4_n_0 ,\fp32_add/Q[87]_i_5_n_0 ,\fp32_add/Q[87]_i_6_n_0 ,\fp32_add/Q[87]_i_7_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[87]_i_3 
       (.CI(\Q_reg[83]_i_3_n_0 ),
        .CO({\Q_reg[87]_i_3_n_1 ,\Q_reg[87]_i_3_n_2 ,\Q_reg[87]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/significand_sub_complement [23:20]),
        .S({\Q[87]_i_8_n_0 ,\Q[87]_i_9_n_0 ,\Q[87]_i_10_n_0 ,\Q[87]_i_11_n_0 }));
  CARRY4 \Q_reg[88]_i_2 
       (.CI(\Q_reg[87]_i_2_n_0 ),
        .CO(\custom_alu/fp32_add/significand_sub0 [24]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \Q_reg[8]_i_1 
       (.CI(\Q_reg[4]_i_1_n_0 ),
        .CO({\Q_reg[8]_i_1_n_0 ,\Q_reg[8]_i_1_n_1 ,\Q_reg[8]_i_1_n_2 ,\Q_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(IF_PC_ADD4[8:5]),
        .S({\Q[8]_i_2__1_n_0 ,\Q[8]_i_3__3_n_0 ,\Q[8]_i_4__2_n_0 ,\Q[8]_i_5__2_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[8]_i_2 
       (.CI(\Q_reg[4]_i_2_n_0 ),
        .CO({\Q_reg[8]_i_2_n_0 ,\Q_reg[8]_i_2_n_1 ,\Q_reg[8]_i_2_n_2 ,\Q_reg[8]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_add/data23 [8:5]),
        .S({\Q[8]_i_4__1_n_0 ,\Q[8]_i_5__0_n_0 ,\Q[8]_i_6__0_n_0 ,\Q[8]_i_7_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[8]_i_2__0 
       (.CI(\Q_reg[4]_i_2__0_n_0 ),
        .CO({\Q_reg[8]_i_2__0_n_0 ,\Q_reg[8]_i_2__0_n_1 ,\Q_reg[8]_i_2__0_n_2 ,\Q_reg[8]_i_2__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/significand_b_add_sub [7:4]),
        .O(\custom_alu/fp32_add/significand_add0 [7:4]),
        .S({\fp32_add/Q[8]_i_7_n_0 ,\fp32_add/Q[8]_i_8_n_0 ,\fp32_add/Q[8]_i_9_n_0 ,\fp32_add/Q[8]_i_10_n_0 }));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \Q_reg[9]_i_5 
       (.CI(\<const0> ),
        .CO({STALL_COUNTER_D1,\Q_reg[9]_i_5_n_1 ,\Q_reg[9]_i_5_n_2 ,\Q_reg[9]_i_5_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\Q[9]_i_8_n_0 ,\Q[9]_i_9__0_n_0 ,\Q[9]_i_10__0_n_0 ,\Q[9]_i_11__0_n_0 }));
  OBUF \RF_RA1_OBUF[0]_inst 
       (.I(CRF_RA1_OBUF[0]),
        .O(RF_RA1[0]));
  OBUF \RF_RA1_OBUF[1]_inst 
       (.I(CRF_RA1_OBUF[1]),
        .O(RF_RA1[1]));
  OBUF \RF_RA1_OBUF[2]_inst 
       (.I(CRF_RA1_OBUF[2]),
        .O(RF_RA1[2]));
  OBUF \RF_RA1_OBUF[3]_inst 
       (.I(CRF_RA1_OBUF[3]),
        .O(RF_RA1[3]));
  OBUF \RF_RA1_OBUF[4]_inst 
       (.I(CRF_RA1_OBUF[4]),
        .O(RF_RA1[4]));
  OBUF \RF_RA2_OBUF[0]_inst 
       (.I(CRF_RA2_OBUF[0]),
        .O(RF_RA2[0]));
  OBUF \RF_RA2_OBUF[1]_inst 
       (.I(CRF_RA2_OBUF[1]),
        .O(RF_RA2[1]));
  OBUF \RF_RA2_OBUF[2]_inst 
       (.I(CRF_RA2_OBUF[2]),
        .O(RF_RA2[2]));
  OBUF \RF_RA2_OBUF[3]_inst 
       (.I(CRF_RA2_OBUF[3]),
        .O(RF_RA2[3]));
  OBUF \RF_RA2_OBUF[4]_inst 
       (.I(CRF_RA2_OBUF[4]),
        .O(RF_RA2[4]));
  IBUF \RF_RD1_IBUF[0]_inst 
       (.I(RF_RD1[0]),
        .O(RF_RD1_IBUF[0]));
  IBUF \RF_RD1_IBUF[10]_inst 
       (.I(RF_RD1[10]),
        .O(RF_RD1_IBUF[10]));
  IBUF \RF_RD1_IBUF[11]_inst 
       (.I(RF_RD1[11]),
        .O(RF_RD1_IBUF[11]));
  IBUF \RF_RD1_IBUF[12]_inst 
       (.I(RF_RD1[12]),
        .O(RF_RD1_IBUF[12]));
  IBUF \RF_RD1_IBUF[13]_inst 
       (.I(RF_RD1[13]),
        .O(RF_RD1_IBUF[13]));
  IBUF \RF_RD1_IBUF[14]_inst 
       (.I(RF_RD1[14]),
        .O(RF_RD1_IBUF[14]));
  IBUF \RF_RD1_IBUF[15]_inst 
       (.I(RF_RD1[15]),
        .O(RF_RD1_IBUF[15]));
  IBUF \RF_RD1_IBUF[16]_inst 
       (.I(RF_RD1[16]),
        .O(RF_RD1_IBUF[16]));
  IBUF \RF_RD1_IBUF[17]_inst 
       (.I(RF_RD1[17]),
        .O(RF_RD1_IBUF[17]));
  IBUF \RF_RD1_IBUF[18]_inst 
       (.I(RF_RD1[18]),
        .O(RF_RD1_IBUF[18]));
  IBUF \RF_RD1_IBUF[19]_inst 
       (.I(RF_RD1[19]),
        .O(RF_RD1_IBUF[19]));
  IBUF \RF_RD1_IBUF[1]_inst 
       (.I(RF_RD1[1]),
        .O(RF_RD1_IBUF[1]));
  IBUF \RF_RD1_IBUF[20]_inst 
       (.I(RF_RD1[20]),
        .O(RF_RD1_IBUF[20]));
  IBUF \RF_RD1_IBUF[21]_inst 
       (.I(RF_RD1[21]),
        .O(RF_RD1_IBUF[21]));
  IBUF \RF_RD1_IBUF[22]_inst 
       (.I(RF_RD1[22]),
        .O(RF_RD1_IBUF[22]));
  IBUF \RF_RD1_IBUF[23]_inst 
       (.I(RF_RD1[23]),
        .O(RF_RD1_IBUF[23]));
  IBUF \RF_RD1_IBUF[24]_inst 
       (.I(RF_RD1[24]),
        .O(RF_RD1_IBUF[24]));
  IBUF \RF_RD1_IBUF[25]_inst 
       (.I(RF_RD1[25]),
        .O(RF_RD1_IBUF[25]));
  IBUF \RF_RD1_IBUF[26]_inst 
       (.I(RF_RD1[26]),
        .O(RF_RD1_IBUF[26]));
  IBUF \RF_RD1_IBUF[27]_inst 
       (.I(RF_RD1[27]),
        .O(RF_RD1_IBUF[27]));
  IBUF \RF_RD1_IBUF[28]_inst 
       (.I(RF_RD1[28]),
        .O(RF_RD1_IBUF[28]));
  IBUF \RF_RD1_IBUF[29]_inst 
       (.I(RF_RD1[29]),
        .O(RF_RD1_IBUF[29]));
  IBUF \RF_RD1_IBUF[2]_inst 
       (.I(RF_RD1[2]),
        .O(RF_RD1_IBUF[2]));
  IBUF \RF_RD1_IBUF[30]_inst 
       (.I(RF_RD1[30]),
        .O(RF_RD1_IBUF[30]));
  IBUF \RF_RD1_IBUF[31]_inst 
       (.I(RF_RD1[31]),
        .O(RF_RD1_IBUF[31]));
  IBUF \RF_RD1_IBUF[3]_inst 
       (.I(RF_RD1[3]),
        .O(RF_RD1_IBUF[3]));
  IBUF \RF_RD1_IBUF[4]_inst 
       (.I(RF_RD1[4]),
        .O(RF_RD1_IBUF[4]));
  IBUF \RF_RD1_IBUF[5]_inst 
       (.I(RF_RD1[5]),
        .O(RF_RD1_IBUF[5]));
  IBUF \RF_RD1_IBUF[6]_inst 
       (.I(RF_RD1[6]),
        .O(RF_RD1_IBUF[6]));
  IBUF \RF_RD1_IBUF[7]_inst 
       (.I(RF_RD1[7]),
        .O(RF_RD1_IBUF[7]));
  IBUF \RF_RD1_IBUF[8]_inst 
       (.I(RF_RD1[8]),
        .O(RF_RD1_IBUF[8]));
  IBUF \RF_RD1_IBUF[9]_inst 
       (.I(RF_RD1[9]),
        .O(RF_RD1_IBUF[9]));
  IBUF \RF_RD2_IBUF[0]_inst 
       (.I(RF_RD2[0]),
        .O(RF_RD2_IBUF[0]));
  IBUF \RF_RD2_IBUF[10]_inst 
       (.I(RF_RD2[10]),
        .O(RF_RD2_IBUF[10]));
  IBUF \RF_RD2_IBUF[11]_inst 
       (.I(RF_RD2[11]),
        .O(RF_RD2_IBUF[11]));
  IBUF \RF_RD2_IBUF[12]_inst 
       (.I(RF_RD2[12]),
        .O(RF_RD2_IBUF[12]));
  IBUF \RF_RD2_IBUF[13]_inst 
       (.I(RF_RD2[13]),
        .O(RF_RD2_IBUF[13]));
  IBUF \RF_RD2_IBUF[14]_inst 
       (.I(RF_RD2[14]),
        .O(RF_RD2_IBUF[14]));
  IBUF \RF_RD2_IBUF[15]_inst 
       (.I(RF_RD2[15]),
        .O(RF_RD2_IBUF[15]));
  IBUF \RF_RD2_IBUF[16]_inst 
       (.I(RF_RD2[16]),
        .O(RF_RD2_IBUF[16]));
  IBUF \RF_RD2_IBUF[17]_inst 
       (.I(RF_RD2[17]),
        .O(RF_RD2_IBUF[17]));
  IBUF \RF_RD2_IBUF[18]_inst 
       (.I(RF_RD2[18]),
        .O(RF_RD2_IBUF[18]));
  IBUF \RF_RD2_IBUF[19]_inst 
       (.I(RF_RD2[19]),
        .O(RF_RD2_IBUF[19]));
  IBUF \RF_RD2_IBUF[1]_inst 
       (.I(RF_RD2[1]),
        .O(RF_RD2_IBUF[1]));
  IBUF \RF_RD2_IBUF[20]_inst 
       (.I(RF_RD2[20]),
        .O(RF_RD2_IBUF[20]));
  IBUF \RF_RD2_IBUF[21]_inst 
       (.I(RF_RD2[21]),
        .O(RF_RD2_IBUF[21]));
  IBUF \RF_RD2_IBUF[22]_inst 
       (.I(RF_RD2[22]),
        .O(RF_RD2_IBUF[22]));
  IBUF \RF_RD2_IBUF[23]_inst 
       (.I(RF_RD2[23]),
        .O(RF_RD2_IBUF[23]));
  IBUF \RF_RD2_IBUF[24]_inst 
       (.I(RF_RD2[24]),
        .O(RF_RD2_IBUF[24]));
  IBUF \RF_RD2_IBUF[25]_inst 
       (.I(RF_RD2[25]),
        .O(RF_RD2_IBUF[25]));
  IBUF \RF_RD2_IBUF[26]_inst 
       (.I(RF_RD2[26]),
        .O(RF_RD2_IBUF[26]));
  IBUF \RF_RD2_IBUF[27]_inst 
       (.I(RF_RD2[27]),
        .O(RF_RD2_IBUF[27]));
  IBUF \RF_RD2_IBUF[28]_inst 
       (.I(RF_RD2[28]),
        .O(RF_RD2_IBUF[28]));
  IBUF \RF_RD2_IBUF[29]_inst 
       (.I(RF_RD2[29]),
        .O(RF_RD2_IBUF[29]));
  IBUF \RF_RD2_IBUF[2]_inst 
       (.I(RF_RD2[2]),
        .O(RF_RD2_IBUF[2]));
  IBUF \RF_RD2_IBUF[30]_inst 
       (.I(RF_RD2[30]),
        .O(RF_RD2_IBUF[30]));
  IBUF \RF_RD2_IBUF[31]_inst 
       (.I(RF_RD2[31]),
        .O(RF_RD2_IBUF[31]));
  IBUF \RF_RD2_IBUF[3]_inst 
       (.I(RF_RD2[3]),
        .O(RF_RD2_IBUF[3]));
  IBUF \RF_RD2_IBUF[4]_inst 
       (.I(RF_RD2[4]),
        .O(RF_RD2_IBUF[4]));
  IBUF \RF_RD2_IBUF[5]_inst 
       (.I(RF_RD2[5]),
        .O(RF_RD2_IBUF[5]));
  IBUF \RF_RD2_IBUF[6]_inst 
       (.I(RF_RD2[6]),
        .O(RF_RD2_IBUF[6]));
  IBUF \RF_RD2_IBUF[7]_inst 
       (.I(RF_RD2[7]),
        .O(RF_RD2_IBUF[7]));
  IBUF \RF_RD2_IBUF[8]_inst 
       (.I(RF_RD2[8]),
        .O(RF_RD2_IBUF[8]));
  IBUF \RF_RD2_IBUF[9]_inst 
       (.I(RF_RD2[9]),
        .O(RF_RD2_IBUF[9]));
  OBUF \RF_WA_OBUF[0]_inst 
       (.I(CRF_WA_OBUF[0]),
        .O(RF_WA[0]));
  OBUF \RF_WA_OBUF[1]_inst 
       (.I(CRF_WA_OBUF[1]),
        .O(RF_WA[1]));
  OBUF \RF_WA_OBUF[2]_inst 
       (.I(CRF_WA_OBUF[2]),
        .O(RF_WA[2]));
  OBUF \RF_WA_OBUF[3]_inst 
       (.I(CRF_WA_OBUF[3]),
        .O(RF_WA[3]));
  OBUF \RF_WA_OBUF[4]_inst 
       (.I(CRF_WA_OBUF[4]),
        .O(RF_WA[4]));
  OBUF \RF_WD_OBUF[0]_inst 
       (.I(CRF_WD_OBUF[0]),
        .O(RF_WD[0]));
  OBUF \RF_WD_OBUF[10]_inst 
       (.I(CRF_WD_OBUF[10]),
        .O(RF_WD[10]));
  OBUF \RF_WD_OBUF[11]_inst 
       (.I(CRF_WD_OBUF[11]),
        .O(RF_WD[11]));
  OBUF \RF_WD_OBUF[12]_inst 
       (.I(CRF_WD_OBUF[12]),
        .O(RF_WD[12]));
  OBUF \RF_WD_OBUF[13]_inst 
       (.I(CRF_WD_OBUF[13]),
        .O(RF_WD[13]));
  OBUF \RF_WD_OBUF[14]_inst 
       (.I(CRF_WD_OBUF[14]),
        .O(RF_WD[14]));
  OBUF \RF_WD_OBUF[15]_inst 
       (.I(CRF_WD_OBUF[15]),
        .O(RF_WD[15]));
  OBUF \RF_WD_OBUF[16]_inst 
       (.I(CRF_WD_OBUF[16]),
        .O(RF_WD[16]));
  OBUF \RF_WD_OBUF[17]_inst 
       (.I(CRF_WD_OBUF[17]),
        .O(RF_WD[17]));
  OBUF \RF_WD_OBUF[18]_inst 
       (.I(CRF_WD_OBUF[18]),
        .O(RF_WD[18]));
  OBUF \RF_WD_OBUF[19]_inst 
       (.I(CRF_WD_OBUF[19]),
        .O(RF_WD[19]));
  OBUF \RF_WD_OBUF[1]_inst 
       (.I(CRF_WD_OBUF[1]),
        .O(RF_WD[1]));
  OBUF \RF_WD_OBUF[20]_inst 
       (.I(CRF_WD_OBUF[20]),
        .O(RF_WD[20]));
  OBUF \RF_WD_OBUF[21]_inst 
       (.I(CRF_WD_OBUF[21]),
        .O(RF_WD[21]));
  OBUF \RF_WD_OBUF[22]_inst 
       (.I(CRF_WD_OBUF[22]),
        .O(RF_WD[22]));
  OBUF \RF_WD_OBUF[23]_inst 
       (.I(CRF_WD_OBUF[23]),
        .O(RF_WD[23]));
  OBUF \RF_WD_OBUF[24]_inst 
       (.I(CRF_WD_OBUF[24]),
        .O(RF_WD[24]));
  OBUF \RF_WD_OBUF[25]_inst 
       (.I(CRF_WD_OBUF[25]),
        .O(RF_WD[25]));
  OBUF \RF_WD_OBUF[26]_inst 
       (.I(CRF_WD_OBUF[26]),
        .O(RF_WD[26]));
  OBUF \RF_WD_OBUF[27]_inst 
       (.I(CRF_WD_OBUF[27]),
        .O(RF_WD[27]));
  OBUF \RF_WD_OBUF[28]_inst 
       (.I(CRF_WD_OBUF[28]),
        .O(RF_WD[28]));
  OBUF \RF_WD_OBUF[29]_inst 
       (.I(CRF_WD_OBUF[29]),
        .O(RF_WD[29]));
  OBUF \RF_WD_OBUF[2]_inst 
       (.I(CRF_WD_OBUF[2]),
        .O(RF_WD[2]));
  OBUF \RF_WD_OBUF[30]_inst 
       (.I(CRF_WD_OBUF[30]),
        .O(RF_WD[30]));
  OBUF \RF_WD_OBUF[31]_inst 
       (.I(CRF_WD_OBUF[31]),
        .O(RF_WD[31]));
  OBUF \RF_WD_OBUF[3]_inst 
       (.I(CRF_WD_OBUF[3]),
        .O(RF_WD[3]));
  OBUF \RF_WD_OBUF[4]_inst 
       (.I(CRF_WD_OBUF[4]),
        .O(RF_WD[4]));
  OBUF \RF_WD_OBUF[5]_inst 
       (.I(CRF_WD_OBUF[5]),
        .O(RF_WD[5]));
  OBUF \RF_WD_OBUF[6]_inst 
       (.I(CRF_WD_OBUF[6]),
        .O(RF_WD[6]));
  OBUF \RF_WD_OBUF[7]_inst 
       (.I(CRF_WD_OBUF[7]),
        .O(RF_WD[7]));
  OBUF \RF_WD_OBUF[8]_inst 
       (.I(CRF_WD_OBUF[8]),
        .O(RF_WD[8]));
  OBUF \RF_WD_OBUF[9]_inst 
       (.I(CRF_WD_OBUF[9]),
        .O(RF_WD[9]));
  OBUF RF_WE_OBUF_inst
       (.I(RF_WE_OBUF),
        .O(RF_WE));
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT2 #(
    .INIT(4'h2)) 
    RF_WE_OBUF_inst_i_1
       (.I0(MEM_WB_Q),
        .I1(WB_CUSTOM_RD),
        .O(RF_WE_OBUF));
  IBUF RSTn_IBUF_inst
       (.I(RSTn),
        .O(RSTn_IBUF));
  VCC VCC
       (.P(\<const1> ));
  VCC VCC_1
       (.P(VCC_2));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [0]),
        .Q(\custom_alu/Q [0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [10]),
        .Q(\custom_alu/Q [10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [11]),
        .Q(\custom_alu/Q [11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [12]),
        .Q(\custom_alu/Q [12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [13]),
        .Q(\custom_alu/Q [13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [14]),
        .Q(\custom_alu/Q [14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [15]),
        .Q(\custom_alu/Q [15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [16]),
        .Q(\custom_alu/Q [16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [17]),
        .Q(\custom_alu/Q [17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [18]),
        .Q(\custom_alu/Q [18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [19]),
        .Q(\custom_alu/Q [19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [1]),
        .Q(\custom_alu/Q [1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [20]),
        .Q(\custom_alu/Q [20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [21]),
        .Q(\custom_alu/Q [21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [22]),
        .Q(\custom_alu/Q [22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [23]),
        .Q(\custom_alu/Q [23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [24]),
        .Q(\custom_alu/Q [24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [25]),
        .Q(\custom_alu/Q [25]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [26]),
        .Q(\custom_alu/Q [26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [27]),
        .Q(\custom_alu/Q [27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [28]),
        .Q(\custom_alu/Q [28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [29]),
        .Q(\custom_alu/Q [29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [2]),
        .Q(\custom_alu/Q [2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [30]),
        .Q(\custom_alu/Q [30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [31]),
        .Q(\custom_alu/Q [31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [3]),
        .Q(\custom_alu/Q [3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [4]),
        .Q(\custom_alu/Q [4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [5]),
        .Q(\custom_alu/Q [5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [6]),
        .Q(\custom_alu/Q [6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [7]),
        .Q(\custom_alu/Q [7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [8]),
        .Q(\custom_alu/Q [8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/FF_FADD/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/FADD_Q [9]),
        .Q(\custom_alu/Q [9]),
        .R(RST0));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp2int/INT0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/fp2int/INT0_carry_n_0 ,\custom_alu/fp2int/INT0_carry_n_1 ,\custom_alu/fp2int/INT0_carry_n_2 ,\custom_alu/fp2int/INT0_carry_n_3 }),
        .CYINIT(\custom_alu/fp2int/p_0_in [0]),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp2int/INT0 [4:1]),
        .S(\custom_alu/fp2int/p_0_in [4:1]));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp2int/INT0_carry__0 
       (.CI(\custom_alu/fp2int/INT0_carry_n_0 ),
        .CO({\custom_alu/fp2int/INT0_carry__0_n_0 ,\custom_alu/fp2int/INT0_carry__0_n_1 ,\custom_alu/fp2int/INT0_carry__0_n_2 ,\custom_alu/fp2int/INT0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp2int/INT0 [8:5]),
        .S(\custom_alu/fp2int/p_0_in [8:5]));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp2int/INT0_carry__1 
       (.CI(\custom_alu/fp2int/INT0_carry__0_n_0 ),
        .CO({\custom_alu/fp2int/INT0_carry__1_n_0 ,\custom_alu/fp2int/INT0_carry__1_n_1 ,\custom_alu/fp2int/INT0_carry__1_n_2 ,\custom_alu/fp2int/INT0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp2int/INT0 [12:9]),
        .S({\custom_alu/fp2int/p_0_in [12],INT0_carry__1_i_2_n_0,\custom_alu/fp2int/p_0_in [10:9]}));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp2int/INT0_carry__2 
       (.CI(\custom_alu/fp2int/INT0_carry__1_n_0 ),
        .CO({\custom_alu/fp2int/INT0_carry__2_n_0 ,\custom_alu/fp2int/INT0_carry__2_n_1 ,\custom_alu/fp2int/INT0_carry__2_n_2 ,\custom_alu/fp2int/INT0_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp2int/INT0 [16:13]),
        .S({INT0_carry__2_i_1_n_0,INT0_carry__2_i_2_n_0,\custom_alu/fp2int/p_0_in [14:13]}));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp2int/INT0_carry__3 
       (.CI(\custom_alu/fp2int/INT0_carry__2_n_0 ),
        .CO({\custom_alu/fp2int/INT0_carry__3_n_0 ,\custom_alu/fp2int/INT0_carry__3_n_1 ,\custom_alu/fp2int/INT0_carry__3_n_2 ,\custom_alu/fp2int/INT0_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp2int/INT0 [20:17]),
        .S({INT0_carry__3_i_1_n_0,INT0_carry__3_i_2_n_0,INT0_carry__3_i_3_n_0,INT0_carry__3_i_4_n_0}));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp2int/INT0_carry__4 
       (.CI(\custom_alu/fp2int/INT0_carry__3_n_0 ),
        .CO({\custom_alu/fp2int/INT0_carry__4_n_0 ,\NLW_custom_alu/fp2int/INT0_carry__4_CO_UNCONNECTED [2],\custom_alu/fp2int/INT0_carry__4_n_2 ,\custom_alu/fp2int/INT0_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp2int/INT0 [23:21]),
        .S({\<const1> ,\custom_alu/fp2int/p_0_in [23],INT0_carry__4_i_2_n_0,\custom_alu/fp2int/p_0_in [21]}));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_in ),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [10]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [11]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [12]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [13]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [14]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [15]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [16]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [17]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [18]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [19]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [1]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [20]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [21]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [22]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [23]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [24]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [25]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [26]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [27]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [28]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [29]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [2]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [30]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [31]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [3]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [4]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [0]),
        .Q(\custom_alu/fp32_add/exp_a [0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [1]),
        .Q(\custom_alu/fp32_add/exp_a [1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [2]),
        .Q(\custom_alu/fp32_add/exp_a [2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [3]),
        .Q(\custom_alu/fp32_add/exp_a [3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [4]),
        .Q(\custom_alu/fp32_add/exp_a [4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [5]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [5]),
        .Q(\custom_alu/fp32_add/exp_a [5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [6]),
        .Q(\custom_alu/fp32_add/exp_a [6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_0_in [7]),
        .Q(\custom_alu/fp32_add/exp_a [7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[64] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [64]),
        .Q(\custom_alu/fp32_add/sel0 [0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[65] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [65]),
        .Q(\custom_alu/fp32_add/sel0 [1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[66] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [66]),
        .Q(\custom_alu/fp32_add/sel0 [2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[67] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [67]),
        .Q(\custom_alu/fp32_add/sel0 [3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[68] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [68]),
        .Q(\custom_alu/fp32_add/sel0 [4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[69] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [69]),
        .Q(\custom_alu/fp32_add/sel0 [5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [6]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[70] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [70]),
        .Q(\custom_alu/fp32_add/sel0 [6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[71] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [71]),
        .Q(\custom_alu/fp32_add/sel0 [7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[72] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [72]),
        .Q(\custom_alu/fp32_add/sel0 [8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[73] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [73]),
        .Q(\custom_alu/fp32_add/sel0 [9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[74] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [74]),
        .Q(\custom_alu/fp32_add/sel0 [10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[75] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [75]),
        .Q(\custom_alu/fp32_add/sel0 [11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[76] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [76]),
        .Q(\custom_alu/fp32_add/sel0 [12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[77] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [77]),
        .Q(\custom_alu/fp32_add/sel0 [13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[78] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [78]),
        .Q(\custom_alu/fp32_add/sel0 [14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[79] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [79]),
        .Q(\custom_alu/fp32_add/sel0 [15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [7]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[80] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [80]),
        .Q(\custom_alu/fp32_add/sel0 [16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[81] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [81]),
        .Q(\custom_alu/fp32_add/sel0 [17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[82] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [82]),
        .Q(\custom_alu/fp32_add/sel0 [18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[83] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [83]),
        .Q(\custom_alu/fp32_add/sel0 [19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[84] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [84]),
        .Q(\custom_alu/fp32_add/sel0 [20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[85] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [85]),
        .Q(\custom_alu/fp32_add/sel0 [21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[86] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [86]),
        .Q(\custom_alu/fp32_add/sel0 [22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[87] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [87]),
        .Q(\custom_alu/fp32_add/sel0 [23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[88] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [88]),
        .Q(\custom_alu/fp32_add/sel0 [24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [8]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_add/FF_PIPELINE/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_add/p_1_out [9]),
        .Q(\custom_alu/fp32_add/FF_PIPELINE/Q_reg_n_0_[9] ),
        .R(RST0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/fp32_add/exp_b_add_sub_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/fp32_add/exp_b_add_sub_carry_n_0 ,\custom_alu/fp32_add/exp_b_add_sub_carry_n_1 ,\custom_alu/fp32_add/exp_b_add_sub_carry_n_2 ,\custom_alu/fp32_add/exp_b_add_sub_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_add/p_0_in2_in [3:0]),
        .O(\custom_alu/fp32_add/exp_b_add_sub [3:0]),
        .S({exp_b_add_sub_carry_i_5_n_0,exp_b_add_sub_carry_i_6_n_0,exp_b_add_sub_carry_i_7_n_0,exp_b_add_sub_carry_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/fp32_add/exp_b_add_sub_carry__0 
       (.CI(\custom_alu/fp32_add/exp_b_add_sub_carry_n_0 ),
        .CO({\custom_alu/fp32_add/exp_b_add_sub_carry__0_n_1 ,\custom_alu/fp32_add/exp_b_add_sub_carry__0_n_2 ,\custom_alu/fp32_add/exp_b_add_sub_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\custom_alu/fp32_add/p_0_in2_in [6:4]}),
        .O(\custom_alu/fp32_add/exp_b_add_sub [7:4]),
        .S({exp_b_add_sub_carry__0_i_4_n_0,exp_b_add_sub_carry__0_i_5_n_0,exp_b_add_sub_carry__0_i_6_n_0,exp_b_add_sub_carry__0_i_7_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/fp32_add/exp_diff_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/fp32_add/exp_diff_carry_n_0 ,\custom_alu/fp32_add/exp_diff_carry_n_1 ,\custom_alu/fp32_add/exp_diff_carry_n_2 ,\custom_alu/fp32_add/exp_diff_carry_n_3 }),
        .CYINIT(\<const1> ),
        .DI({exp_diff_carry_i_1_n_0,exp_diff_carry_i_2_n_0,exp_diff_carry_i_3_n_0,exp_diff_carry_i_4_n_0}),
        .O(\custom_alu/fp32_add/p_1_in__0 [3:0]),
        .S({exp_diff_carry_i_5_n_0,exp_diff_carry_i_6_n_0,exp_diff_carry_i_7_n_0,exp_diff_carry_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/fp32_add/exp_diff_carry__0 
       (.CI(\custom_alu/fp32_add/exp_diff_carry_n_0 ),
        .CO({\custom_alu/fp32_add/exp_diff_carry__0_n_1 ,\custom_alu/fp32_add/exp_diff_carry__0_n_2 ,\custom_alu/fp32_add/exp_diff_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,exp_diff_carry__0_i_1_n_0,exp_diff_carry__0_i_2_n_0,exp_diff_carry__0_i_3_n_0}),
        .O(\custom_alu/fp32_add/p_1_in__0 [7:4]),
        .S({exp_diff_carry__0_i_4_n_0,exp_diff_carry__0_i_5_n_0,exp_diff_carry__0_i_6_n_0,exp_diff_carry__0_i_7_n_0}));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \custom_alu/fp32_add/op_a2_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/fp32_add/op_a2_carry_n_0 ,\custom_alu/fp32_add/op_a2_carry_n_1 ,\custom_alu/fp32_add/op_a2_carry_n_2 ,\custom_alu/fp32_add/op_a2_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({op_a2_carry_i_1_n_0,op_a2_carry_i_2_n_0,op_a2_carry_i_3_n_0,op_a2_carry_i_4_n_0}),
        .S({op_a2_carry_i_5_n_0,op_a2_carry_i_6_n_0,op_a2_carry_i_7_n_0,op_a2_carry_i_8_n_0}));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \custom_alu/fp32_add/op_a2_carry__0 
       (.CI(\custom_alu/fp32_add/op_a2_carry_n_0 ),
        .CO({\custom_alu/fp32_add/op_a2_carry__0_n_0 ,\custom_alu/fp32_add/op_a2_carry__0_n_1 ,\custom_alu/fp32_add/op_a2_carry__0_n_2 ,\custom_alu/fp32_add/op_a2_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({op_a2_carry__0_i_1_n_0,op_a2_carry__0_i_2_n_0,op_a2_carry__0_i_3_n_0,op_a2_carry__0_i_4_n_0}),
        .S({op_a2_carry__0_i_5_n_0,op_a2_carry__0_i_6_n_0,op_a2_carry__0_i_7_n_0,op_a2_carry__0_i_8_n_0}));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \custom_alu/fp32_add/op_a2_carry__1 
       (.CI(\custom_alu/fp32_add/op_a2_carry__0_n_0 ),
        .CO({\custom_alu/fp32_add/op_a2_carry__1_n_0 ,\custom_alu/fp32_add/op_a2_carry__1_n_1 ,\custom_alu/fp32_add/op_a2_carry__1_n_2 ,\custom_alu/fp32_add/op_a2_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({op_a2_carry__1_i_1_n_0,op_a2_carry__1_i_2_n_0,op_a2_carry__1_i_3_n_0,op_a2_carry__1_i_4_n_0}),
        .S({op_a2_carry__1_i_5_n_0,op_a2_carry__1_i_6_n_0,op_a2_carry__1_i_7_n_0,op_a2_carry__1_i_8_n_0}));
  (* COMPARATOR_THRESHOLD = "11" *) 
  CARRY4 \custom_alu/fp32_add/op_a2_carry__2 
       (.CI(\custom_alu/fp32_add/op_a2_carry__1_n_0 ),
        .CO({\custom_alu/fp32_add/op_a2 ,\custom_alu/fp32_add/op_a2_carry__2_n_1 ,\custom_alu/fp32_add/op_a2_carry__2_n_2 ,\custom_alu/fp32_add/op_a2_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({op_a2_carry__2_i_1_n_0,op_a2_carry__2_i_2_n_0,op_a2_carry__2_i_3_n_0,op_a2_carry__2_i_4_n_0}),
        .S({op_a2_carry__2_i_5_n_0,op_a2_carry__2_i_6_n_0,op_a2_carry__2_i_7_n_0,op_a2_carry__2_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp32_add/pe/exp_sub_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/fp32_add/pe/exp_sub_carry_n_0 ,\custom_alu/fp32_add/pe/exp_sub_carry_n_1 ,\custom_alu/fp32_add/pe/exp_sub_carry_n_2 ,\custom_alu/fp32_add/pe/exp_sub_carry_n_3 }),
        .CYINIT(\<const1> ),
        .DI(\custom_alu/fp32_add/exp_a [3:0]),
        .O(\custom_alu/fp32_add/exp_sub [3:0]),
        .S({exp_sub_carry_i_1_n_0,exp_sub_carry_i_2_n_0,exp_sub_carry_i_3_n_0,exp_sub_carry_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp32_add/pe/exp_sub_carry__0 
       (.CI(\custom_alu/fp32_add/pe/exp_sub_carry_n_0 ),
        .CO({\custom_alu/fp32_add/pe/exp_sub_carry__0_n_1 ,\custom_alu/fp32_add/pe/exp_sub_carry__0_n_2 ,\custom_alu/fp32_add/pe/exp_sub_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\custom_alu/fp32_add/exp_a [6:4]}),
        .O(\custom_alu/fp32_add/exp_sub [7:4]),
        .S({exp_sub_carry__0_i_1_n_0,exp_sub_carry__0_i_2_n_0,exp_sub_carry__0_i_3_n_0,exp_sub_carry__0_i_4_n_0}));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[23]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[24]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[25]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[26]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[27]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[28]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[29]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[30]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN2[31]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[23]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[24]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[25]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[26]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[27]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[28]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[29]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(ALU_DIN1[30]),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_1/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\Q[63]_i_1__1_n_0 ),
        .Q(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[63] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[23] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[24] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[25] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[26] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[27] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[28] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[29] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[30] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[31] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[55] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[56] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[57] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[58] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[59] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[60] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[61] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[62] ),
        .Q(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/FF_MULT_2/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/FF_MULT_1/Q_reg_n_0_[63] ),
        .Q(\custom_alu/fp32_mult/a_Q ),
        .R(RST0));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp32_mult/exponent_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/fp32_mult/exponent_carry_n_0 ,\custom_alu/fp32_mult/exponent_carry_n_1 ,\custom_alu/fp32_mult/exponent_carry_n_2 ,\custom_alu/fp32_mult/exponent_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({exponent_carry_i_1_n_0,exponent_carry_i_2_n_0,exponent_carry_i_3_n_0,\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[55] }),
        .O({\custom_alu/fp32_mult/exponent_carry_n_4 ,\custom_alu/fp32_mult/exponent_carry_n_5 ,\custom_alu/fp32_mult/exponent_carry_n_6 ,\custom_alu/fp32_mult/exponent_carry_n_7 }),
        .S({exponent_carry_i_4_n_0,exponent_carry_i_5_n_0,exponent_carry_i_6_n_0,exponent_carry_i_7_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp32_mult/exponent_carry__0 
       (.CI(\custom_alu/fp32_mult/exponent_carry_n_0 ),
        .CO({\custom_alu/fp32_mult/exponent_carry__0_n_0 ,\custom_alu/fp32_mult/exponent_carry__0_n_1 ,\custom_alu/fp32_mult/exponent_carry__0_n_2 ,\custom_alu/fp32_mult/exponent_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({exponent_carry__0_i_1_n_0,exponent_carry__0_i_2_n_0,exponent_carry__0_i_3_n_0,exponent_carry__0_i_4_n_0}),
        .O({\custom_alu/fp32_mult/p_0_in1_in ,\custom_alu/fp32_mult/exponent_carry__0_n_5 ,\custom_alu/fp32_mult/exponent_carry__0_n_6 ,\custom_alu/fp32_mult/exponent_carry__0_n_7 }),
        .S({exponent_carry__0_i_5_n_0,exponent_carry__0_i_6_n_0,exponent_carry__0_i_7_n_0,exponent_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \custom_alu/fp32_mult/exponent_carry__1 
       (.CI(\custom_alu/fp32_mult/exponent_carry__0_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_mult/exponent_carry__1_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,exponent_carry__1_i_1_n_0}));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [0]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [10]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [11]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [12]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [13]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [14]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [15]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [16]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [17]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [18]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [19]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [1]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [20]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [21]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [22]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [23]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [24]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [0]),
        .Q(\custom_alu/fp32_mult/p_1_in [0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [1]),
        .Q(\custom_alu/fp32_mult/p_1_in [1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [2]),
        .Q(\custom_alu/fp32_mult/p_1_in [2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [3]),
        .Q(\custom_alu/fp32_mult/p_1_in [3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [4]),
        .Q(\custom_alu/fp32_mult/p_1_in [4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [2]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [5]),
        .Q(\custom_alu/fp32_mult/p_1_in [5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [6]),
        .Q(\custom_alu/fp32_mult/p_1_in [6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [7]),
        .Q(\custom_alu/fp32_mult/p_1_in [7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [8]),
        .Q(\custom_alu/fp32_mult/p_1_in [8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [9]),
        .Q(\custom_alu/fp32_mult/p_1_in [9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [10]),
        .Q(\custom_alu/fp32_mult/p_1_in [10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [11]),
        .Q(\custom_alu/fp32_mult/p_1_in [11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [12]),
        .Q(\custom_alu/fp32_mult/p_1_in [12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [13]),
        .Q(\custom_alu/fp32_mult/p_1_in [13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [14]),
        .Q(\custom_alu/fp32_mult/p_1_in [14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [3]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [15]),
        .Q(\custom_alu/fp32_mult/p_1_in [15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [16]),
        .Q(\custom_alu/fp32_mult/p_1_in [16]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [17]),
        .Q(\custom_alu/fp32_mult/p_1_in [17]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [18]),
        .Q(\custom_alu/fp32_mult/p_1_in [18]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [19]),
        .Q(\custom_alu/fp32_mult/p_1_in [19]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [20]),
        .Q(\custom_alu/fp32_mult/p_1_in [20]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [21]),
        .Q(\custom_alu/fp32_mult/p_1_in [21]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [22]),
        .Q(\custom_alu/fp32_mult/p_1_in [22]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM0__0 [23]),
        .Q(\custom_alu/fp32_mult/p_1_in [23]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[49] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [0]),
        .Q(\custom_alu/fp32_mult/p_1_in [24]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [4]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[50] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [1]),
        .Q(\custom_alu/fp32_mult/p_1_in [25]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[51] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [2]),
        .Q(\custom_alu/fp32_mult/p_1_in [26]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[52] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [3]),
        .Q(\custom_alu/fp32_mult/p_1_in [27]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[53] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [4]),
        .Q(\custom_alu/fp32_mult/p_1_in [28]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[54] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [5]),
        .Q(\custom_alu/fp32_mult/p_1_in [29]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [6]),
        .Q(\custom_alu/fp32_mult/p_1_in [30]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [7]),
        .Q(\custom_alu/fp32_mult/p_1_in [31]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [8]),
        .Q(\custom_alu/fp32_mult/p_1_in [32]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [9]),
        .Q(\custom_alu/fp32_mult/p_1_in [33]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [10]),
        .Q(\custom_alu/fp32_mult/p_1_in [34]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [5]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [11]),
        .Q(\custom_alu/fp32_mult/p_1_in [35]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [12]),
        .Q(\custom_alu/fp32_mult/p_1_in [36]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [13]),
        .Q(\custom_alu/fp32_mult/p_1_in [37]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [14]),
        .Q(\custom_alu/fp32_mult/p_1_in [38]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[64] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [15]),
        .Q(\custom_alu/fp32_mult/p_1_in [39]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[65] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [16]),
        .Q(\custom_alu/fp32_mult/p_1_in [40]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[66] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [17]),
        .Q(\custom_alu/fp32_mult/p_1_in [41]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[67] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [18]),
        .Q(\custom_alu/fp32_mult/p_1_in [42]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[68] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [19]),
        .Q(\custom_alu/fp32_mult/p_1_in [43]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[69] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [20]),
        .Q(\custom_alu/fp32_mult/p_1_in [44]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [6]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[70] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [21]),
        .Q(\custom_alu/fp32_mult/p_1_in [45]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[71] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [22]),
        .Q(\custom_alu/fp32_mult/p_1_in [46]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[72] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/mult24_0/PSUM3__0 [23]),
        .Q(\custom_alu/fp32_mult/p_1_in [47]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [7]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [8]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/fp32_mult/PSUM1_2 [9]),
        .Q(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[9] ),
        .R(RST0));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \custom_alu/fp32_mult/mult24_0/PSUM0 
       (.A({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,ALU_DIN1[11:0]}),
        .ACIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .ALUMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .B({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,ALU_DIN2[11:0]}),
        .BCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0> ),
        .CARRYIN(\<const0> ),
        .CARRYINSEL({\<const0> ,\<const0> ,\<const0> }),
        .CEA1(\<const0> ),
        .CEA2(\<const0> ),
        .CEAD(\<const0> ),
        .CEALUMODE(\<const0> ),
        .CEB1(\<const0> ),
        .CEB2(\<const0> ),
        .CEC(\<const0> ),
        .CECARRYIN(\<const0> ),
        .CECTRL(\<const0> ),
        .CED(\<const0> ),
        .CEINMODE(\<const0> ),
        .CEM(\<const0> ),
        .CEP(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .MULTSIGNIN(\<const0> ),
        .OPMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const1> ,\<const0> ,\<const1> }),
        .P(\custom_alu/fp32_mult/mult24_0/PSUM0__0 ),
        .PCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .RSTA(\<const0> ),
        .RSTALLCARRYIN(\<const0> ),
        .RSTALUMODE(\<const0> ),
        .RSTB(\<const0> ),
        .RSTC(\<const0> ),
        .RSTCTRL(\<const0> ),
        .RSTD(\<const0> ),
        .RSTINMODE(\<const0> ),
        .RSTM(\<const0> ),
        .RSTP(RST0));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \custom_alu/fp32_mult/mult24_0/PSUM1 
       (.A({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\custom_alu/fp32_mult/op_a1 ,ALU_DIN1[22:12]}),
        .ACIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .ALUMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .B({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,ALU_DIN2[11:0]}),
        .BCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0> ),
        .CARRYIN(\<const0> ),
        .CARRYINSEL({\<const0> ,\<const0> ,\<const0> }),
        .CEA1(\<const0> ),
        .CEA2(\<const0> ),
        .CEAD(\<const0> ),
        .CEALUMODE(\<const0> ),
        .CEB1(\<const0> ),
        .CEB2(\<const0> ),
        .CEC(\<const0> ),
        .CECARRYIN(\<const0> ),
        .CECTRL(\<const0> ),
        .CED(\<const0> ),
        .CEINMODE(\<const0> ),
        .CEM(\<const0> ),
        .CEP(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .MULTSIGNIN(\<const0> ),
        .OPMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const1> ,\<const0> ,\<const1> }),
        .P(\custom_alu/fp32_mult/mult24_0/PSUM1__0 ),
        .PCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .RSTA(\<const0> ),
        .RSTALLCARRYIN(\<const0> ),
        .RSTALUMODE(\<const0> ),
        .RSTB(\<const0> ),
        .RSTC(\<const0> ),
        .RSTCTRL(\<const0> ),
        .RSTD(\<const0> ),
        .RSTINMODE(\<const0> ),
        .RSTM(\<const0> ),
        .RSTP(RST0));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \custom_alu/fp32_mult/mult24_0/PSUM2 
       (.A({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,ALU_DIN1[11:0]}),
        .ACIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .ALUMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .B({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\custom_alu/fp32_mult/op_b1 ,ALU_DIN2[22:12]}),
        .BCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0> ),
        .CARRYIN(\<const0> ),
        .CARRYINSEL({\<const0> ,\<const0> ,\<const0> }),
        .CEA1(\<const0> ),
        .CEA2(\<const0> ),
        .CEAD(\<const0> ),
        .CEALUMODE(\<const0> ),
        .CEB1(\<const0> ),
        .CEB2(\<const0> ),
        .CEC(\<const0> ),
        .CECARRYIN(\<const0> ),
        .CECTRL(\<const0> ),
        .CED(\<const0> ),
        .CEINMODE(\<const0> ),
        .CEM(\<const0> ),
        .CEP(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .MULTSIGNIN(\<const0> ),
        .OPMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const1> ,\<const0> ,\<const1> }),
        .P(\custom_alu/fp32_mult/p_0_in ),
        .PCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .RSTA(\<const0> ),
        .RSTALLCARRYIN(\<const0> ),
        .RSTALUMODE(\<const0> ),
        .RSTB(\<const0> ),
        .RSTC(\<const0> ),
        .RSTCTRL(\<const0> ),
        .RSTD(\<const0> ),
        .RSTINMODE(\<const0> ),
        .RSTM(\<const0> ),
        .RSTP(RST0));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \custom_alu/fp32_mult/mult24_0/PSUM3 
       (.A({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\custom_alu/fp32_mult/op_a1 ,ALU_DIN1[22:12]}),
        .ACIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .ALUMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .B({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\custom_alu/fp32_mult/op_b1 ,ALU_DIN2[22:12]}),
        .BCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0> ),
        .CARRYIN(\<const0> ),
        .CARRYINSEL({\<const0> ,\<const0> ,\<const0> }),
        .CEA1(\<const0> ),
        .CEA2(\<const0> ),
        .CEAD(\<const0> ),
        .CEALUMODE(\<const0> ),
        .CEB1(\<const0> ),
        .CEB2(\<const0> ),
        .CEC(\<const0> ),
        .CECARRYIN(\<const0> ),
        .CECTRL(\<const0> ),
        .CED(\<const0> ),
        .CEINMODE(\<const0> ),
        .CEM(\<const0> ),
        .CEP(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .MULTSIGNIN(\<const0> ),
        .OPMODE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const1> ,\<const0> ,\<const1> }),
        .P(\custom_alu/fp32_mult/mult24_0/PSUM3__0 ),
        .PCIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .RSTA(\<const0> ),
        .RSTALLCARRYIN(\<const0> ),
        .RSTALUMODE(\<const0> ),
        .RSTB(\<const0> ),
        .RSTC(\<const0> ),
        .RSTCTRL(\<const0> ),
        .RSTD(\<const0> ),
        .RSTINMODE(\<const0> ),
        .RSTM(\<const0> ),
        .RSTP(RST0));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[11]_i_2 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [11]),
        .I1(\custom_alu/fp32_mult/p_0_in [11]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[11]_i_3 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [10]),
        .I1(\custom_alu/fp32_mult/p_0_in [10]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[11]_i_4 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [9]),
        .I1(\custom_alu/fp32_mult/p_0_in [9]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[11]_i_5 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [8]),
        .I1(\custom_alu/fp32_mult/p_0_in [8]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[15]_i_2 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [15]),
        .I1(\custom_alu/fp32_mult/p_0_in [15]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[15]_i_3 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [14]),
        .I1(\custom_alu/fp32_mult/p_0_in [14]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[15]_i_4 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [13]),
        .I1(\custom_alu/fp32_mult/p_0_in [13]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[15]_i_5 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [12]),
        .I1(\custom_alu/fp32_mult/p_0_in [12]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[19]_i_2 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [19]),
        .I1(\custom_alu/fp32_mult/p_0_in [19]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[19]_i_3 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [18]),
        .I1(\custom_alu/fp32_mult/p_0_in [18]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[19]_i_4 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [17]),
        .I1(\custom_alu/fp32_mult/p_0_in [17]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[19]_i_5 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [16]),
        .I1(\custom_alu/fp32_mult/p_0_in [16]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[19]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[23]_i_2 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [23]),
        .I1(\custom_alu/fp32_mult/p_0_in [23]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[23]_i_3 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [22]),
        .I1(\custom_alu/fp32_mult/p_0_in [22]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[23]_i_4 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [21]),
        .I1(\custom_alu/fp32_mult/p_0_in [21]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[23]_i_5 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [20]),
        .I1(\custom_alu/fp32_mult/p_0_in [20]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[23]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[3]_i_2 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [3]),
        .I1(\custom_alu/fp32_mult/p_0_in [3]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[3]_i_3 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [2]),
        .I1(\custom_alu/fp32_mult/p_0_in [2]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[3]_i_4 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [1]),
        .I1(\custom_alu/fp32_mult/p_0_in [1]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[3]_i_5 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [0]),
        .I1(\custom_alu/fp32_mult/p_0_in [0]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[7]_i_2 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [7]),
        .I1(\custom_alu/fp32_mult/p_0_in [7]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[7]_i_3 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [6]),
        .I1(\custom_alu/fp32_mult/p_0_in [6]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[7]_i_4 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [5]),
        .I1(\custom_alu/fp32_mult/p_0_in [5]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/fp32_mult/mult24_0/Q[7]_i_5 
       (.I0(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [4]),
        .I1(\custom_alu/fp32_mult/p_0_in [4]),
        .O(\custom_alu/fp32_mult/mult24_0/Q[7]_i_5_n_0 ));
  CARRY4 \custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1 
       (.CI(\custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_0 ),
        .CO({\custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_0 ,\custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_1 ,\custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_2 ,\custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [11:8]),
        .O(\custom_alu/fp32_mult/PSUM1_2 [11:8]),
        .S({\custom_alu/fp32_mult/mult24_0/Q[11]_i_2_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[11]_i_3_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[11]_i_4_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[11]_i_5_n_0 }));
  CARRY4 \custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1 
       (.CI(\custom_alu/fp32_mult/mult24_0/Q_reg[11]_i_1_n_0 ),
        .CO({\custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_0 ,\custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_1 ,\custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_2 ,\custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [15:12]),
        .O(\custom_alu/fp32_mult/PSUM1_2 [15:12]),
        .S({\custom_alu/fp32_mult/mult24_0/Q[15]_i_2_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[15]_i_3_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[15]_i_4_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[15]_i_5_n_0 }));
  CARRY4 \custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1 
       (.CI(\custom_alu/fp32_mult/mult24_0/Q_reg[15]_i_1_n_0 ),
        .CO({\custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_0 ,\custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_1 ,\custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_2 ,\custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [19:16]),
        .O(\custom_alu/fp32_mult/PSUM1_2 [19:16]),
        .S({\custom_alu/fp32_mult/mult24_0/Q[19]_i_2_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[19]_i_3_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[19]_i_4_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[19]_i_5_n_0 }));
  CARRY4 \custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1 
       (.CI(\custom_alu/fp32_mult/mult24_0/Q_reg[19]_i_1_n_0 ),
        .CO({\custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_0 ,\custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_1 ,\custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_2 ,\custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [23:20]),
        .O(\custom_alu/fp32_mult/PSUM1_2 [23:20]),
        .S({\custom_alu/fp32_mult/mult24_0/Q[23]_i_2_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[23]_i_3_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[23]_i_4_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[23]_i_5_n_0 }));
  CARRY4 \custom_alu/fp32_mult/mult24_0/Q_reg[24]_i_1 
       (.CI(\custom_alu/fp32_mult/mult24_0/Q_reg[23]_i_1_n_0 ),
        .CO(\custom_alu/fp32_mult/PSUM1_2 [24]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  CARRY4 \custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_0 ,\custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_1 ,\custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_2 ,\custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [3:0]),
        .O(\custom_alu/fp32_mult/PSUM1_2 [3:0]),
        .S({\custom_alu/fp32_mult/mult24_0/Q[3]_i_2_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[3]_i_3_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[3]_i_4_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[3]_i_5_n_0 }));
  CARRY4 \custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1 
       (.CI(\custom_alu/fp32_mult/mult24_0/Q_reg[3]_i_1_n_0 ),
        .CO({\custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_0 ,\custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_1 ,\custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_2 ,\custom_alu/fp32_mult/mult24_0/Q_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/fp32_mult/mult24_0/PSUM1__0 [7:4]),
        .O(\custom_alu/fp32_mult/PSUM1_2 [7:4]),
        .S({\custom_alu/fp32_mult/mult24_0/Q[7]_i_2_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[7]_i_3_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[7]_i_4_n_0 ,\custom_alu/fp32_mult/mult24_0/Q[7]_i_5_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[0]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[0]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[100]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[100]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[101]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[101]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[102]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[102]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[103] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [7]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[103] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[104] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [8]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[104] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[105] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [9]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[105] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[106] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [10]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[106] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[107] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [11]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[107] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[108] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [12]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[108] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[109] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [13]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[109] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[110] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [14]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[110] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[111] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [15]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[111] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[112] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [16]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[112] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[113] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [17]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[113] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[114] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [18]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[114] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[115] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [19]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[115] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[116] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [20]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[116] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[117] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [21]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[117] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[118] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [22]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[118] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[119] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [23]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[119] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[120] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [24]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[120] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[121] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [25]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[121] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[122] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [26]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[122] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[123] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [27]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[123] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[124] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [28]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[124] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[125] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [29]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[125] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[126] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [30]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[126] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[127] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0_1_2_3 [31]),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[127] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[1]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[1]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[2]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[2]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[31]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[17] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[18] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[19] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[20] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[21] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[22] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[23] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[3]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[3]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[49] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[49] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[4]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[4]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[50] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[50] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[51] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[51] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[52] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[52] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[53] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[53] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[54] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[54] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[5]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[5]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[63]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[63] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[64] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[17] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[64] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[65] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[18] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[65] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[66] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[19] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[66] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[67] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[20] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[67] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[68] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[21] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[68] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[69] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[22] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[69] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[6]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[6]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[70] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[23] ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[70] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[71] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[71] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[72] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[72] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[73] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[73] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[74] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[74] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[75] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[75] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[76] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[76] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[77] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[77] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[78] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[78] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[79] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[79] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[80] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[80] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[81] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[81] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[82] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[82] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[83] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[83] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[84] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[84] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[85] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[85] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[86] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[86] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[87] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[87] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[88] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[88] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[89] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[89] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[90] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[90] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[91] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[91] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[92] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[92] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[93] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[93] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[94] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[94] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[95] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[95]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[95] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[96]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[96]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[97]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[97]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[98]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[98]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[99]_custom_alu_mult_FF_MULT_0_Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg[99]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[9] ),
        .R(RST0));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[6]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__0 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[5]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__0_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__1 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[4]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__10 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[98]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__10_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__11 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[97]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__11_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__12 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[96]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__12_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[3]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[2]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[1]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[0]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__5_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__6 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[102]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__6_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__7 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[101]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__7_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__8 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[100]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__8_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_gate__9 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg[99]_custom_alu_mult_FF_MULT_0_Q_reg_r_n_0 ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .O(\custom_alu/mult/FF_MULT_0/Q_reg_gate__9_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_0/Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_0/Q_reg_r_n_0 ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[3]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[11]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[11]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[15]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[15]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[15]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[15]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[19]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[19]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[19]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[19]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[3]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[23]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[23]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[23]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[23]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[27]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[27]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[27]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[27]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[31]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[31]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[3]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[31]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[31]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[32]_i_1_n_3 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__12_n_0 ),
        .Q(\custom_alu/MULT [0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__11_n_0 ),
        .Q(\custom_alu/MULT [1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__10_n_0 ),
        .Q(\custom_alu/MULT [2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__9_n_0 ),
        .Q(\custom_alu/MULT [3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__8_n_0 ),
        .Q(\custom_alu/MULT [4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__7_n_0 ),
        .Q(\custom_alu/MULT [5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__6_n_0 ),
        .Q(\custom_alu/MULT [6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[3]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[103] ),
        .Q(\custom_alu/MULT [7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[104] ),
        .Q(\custom_alu/MULT [8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[105] ),
        .Q(\custom_alu/MULT [9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[106] ),
        .Q(\custom_alu/MULT [10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[107] ),
        .Q(\custom_alu/MULT [11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[108] ),
        .Q(\custom_alu/MULT [12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[109] ),
        .Q(\custom_alu/MULT [13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[110] ),
        .Q(\custom_alu/MULT [14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[111] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[49] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[112] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[49] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[7]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[50] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[113] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[50] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[51] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[114] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[51] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[52] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[115] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[52] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[53] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[116] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[53] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[54] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[117] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[54] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[118] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[119] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[120] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[121] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[122] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[7]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[123] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[124] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[125] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[126] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[63] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[64] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[127] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[64] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[65] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__5_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[65] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[66] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__4_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[66] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[67] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__3_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[67] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[68] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__2_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[68] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[69] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__1_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[69] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[7]_i_1_n_5 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[70] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate__0_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[70] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[71] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_gate_n_0 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[71] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[72] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[7] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[72] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[73] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[8] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[73] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[74] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[9] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[74] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[75] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[10] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[75] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[76] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[11] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[76] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[77] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[12] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[77] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[78] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[13] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[78] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[79] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[14] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[79] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[7]_i_1_n_4 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[80] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[15] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[80] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[81] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[16] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[81] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[82] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[17] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[82] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[83] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[18] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[83] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[84] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[19] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[84] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[85] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[20] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[85] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[86] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[21] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[86] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[87] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[22] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[87] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[88] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[23] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[88] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[89] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[24] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[89] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[11]_i_1_n_7 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[90] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[25] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[90] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[91] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[26] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[91] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[92] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[27] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[92] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[93] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[28] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[93] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[94] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[29] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[94] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[95] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[30] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[95] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[96] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[31] ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[96] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/FF_MULT_1/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/Q_reg[11]_i_1_n_6 ),
        .Q(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[9] ),
        .R(RST0));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_12 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[71] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[22] ),
        .O(\custom_alu/mult/Q[11]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_13 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[70] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[21] ),
        .O(\custom_alu/mult/Q[11]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_14 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[69] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[20] ),
        .O(\custom_alu/mult/Q[11]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_15 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[68] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[19] ),
        .O(\custom_alu/mult/Q[11]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[43] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[75] ),
        .O(\custom_alu/mult/Q[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[42] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[74] ),
        .O(\custom_alu/mult/Q[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[73] ),
        .O(\custom_alu/mult/Q[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[11]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[72] ),
        .O(\custom_alu/mult/Q[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_10 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[73] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[24] ),
        .O(\custom_alu/mult/Q[15]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_11 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[72] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[23] ),
        .O(\custom_alu/mult/Q[15]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[47] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[79] ),
        .O(\custom_alu/mult/Q[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[46] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[78] ),
        .O(\custom_alu/mult/Q[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[45] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[77] ),
        .O(\custom_alu/mult/Q[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[44] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[76] ),
        .O(\custom_alu/mult/Q[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_8 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[75] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[26] ),
        .O(\custom_alu/mult/Q[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[15]_i_9 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[74] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[25] ),
        .O(\custom_alu/mult/Q[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_10 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[77] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[28] ),
        .O(\custom_alu/mult/Q[19]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_11 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[76] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[27] ),
        .O(\custom_alu/mult/Q[19]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[51] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[83] ),
        .O(\custom_alu/mult/Q[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[50] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[82] ),
        .O(\custom_alu/mult/Q[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[49] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[81] ),
        .O(\custom_alu/mult/Q[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[48] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[80] ),
        .O(\custom_alu/mult/Q[19]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_8 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[79] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[30] ),
        .O(\custom_alu/mult/Q[19]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[19]_i_9 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[78] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[29] ),
        .O(\custom_alu/mult/Q[19]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_10 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[49] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[0] ),
        .O(\custom_alu/mult/Q[23]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_11 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[81] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[32] ),
        .O(\custom_alu/mult/Q[23]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_12 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[80] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[31] ),
        .O(\custom_alu/mult/Q[23]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[55] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[87] ),
        .O(\custom_alu/mult/Q[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[54] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[86] ),
        .O(\custom_alu/mult/Q[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[53] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[85] ),
        .O(\custom_alu/mult/Q[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[52] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[84] ),
        .O(\custom_alu/mult/Q[23]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_8 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[51] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[2] ),
        .O(\custom_alu/mult/Q[23]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[23]_i_9 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[50] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[1] ),
        .O(\custom_alu/mult/Q[23]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_10 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[54] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[5] ),
        .O(\custom_alu/mult/Q[27]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_11 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[53] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[4] ),
        .O(\custom_alu/mult/Q[27]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_12 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[52] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[3] ),
        .O(\custom_alu/mult/Q[27]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[59] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[91] ),
        .O(\custom_alu/mult/Q[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[58] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[90] ),
        .O(\custom_alu/mult/Q[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[57] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[89] ),
        .O(\custom_alu/mult/Q[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[56] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[88] ),
        .O(\custom_alu/mult/Q[27]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[27]_i_9 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[55] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[6] ),
        .O(\custom_alu/mult/Q[27]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_15 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[59] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[10] ),
        .O(\custom_alu/mult/Q[31]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_16 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[58] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[9] ),
        .O(\custom_alu/mult/Q[31]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_17 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[57] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[8] ),
        .O(\custom_alu/mult/Q[31]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_18 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[56] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[7] ),
        .O(\custom_alu/mult/Q[31]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[63] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[95] ),
        .O(\custom_alu/mult/Q[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[62] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[94] ),
        .O(\custom_alu/mult/Q[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[61] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[93] ),
        .O(\custom_alu/mult/Q[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[31]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[60] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[92] ),
        .O(\custom_alu/mult/Q[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[35]_i_12 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[63] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[14] ),
        .O(\custom_alu/mult/Q[35]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[35]_i_13 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[62] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[13] ),
        .O(\custom_alu/mult/Q[35]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[35]_i_14 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[61] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[12] ),
        .O(\custom_alu/mult/Q[35]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[35]_i_15 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[60] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[11] ),
        .O(\custom_alu/mult/Q[35]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[3]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[67] ),
        .O(\custom_alu/mult/Q[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[3]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[66] ),
        .O(\custom_alu/mult/Q[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[3]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[65] ),
        .O(\custom_alu/mult/Q[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[3]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[64] ),
        .O(\custom_alu/mult/Q[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[5]_i_6 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[67] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[18] ),
        .O(\custom_alu/mult/Q[5]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[5]_i_7 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[66] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[17] ),
        .O(\custom_alu/mult/Q[5]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[5]_i_8 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[65] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/Q[5]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[5]_i_9 
       (.I0(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[64] ),
        .I1(\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[15] ),
        .O(\custom_alu/mult/Q[5]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[7]_i_2 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[71] ),
        .O(\custom_alu/mult/Q[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[7]_i_3 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[70] ),
        .O(\custom_alu/mult/Q[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[7]_i_4 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[69] ),
        .O(\custom_alu/mult/Q[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/Q[7]_i_5 
       (.I0(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[68] ),
        .O(\custom_alu/mult/Q[7]_i_5_n_0 ));
  CARRY4 \custom_alu/mult/Q_reg[11]_i_1 
       (.CI(\custom_alu/mult/Q_reg[7]_i_1_n_0 ),
        .CO({\custom_alu/mult/Q_reg[11]_i_1_n_0 ,\custom_alu/mult/Q_reg[11]_i_1_n_1 ,\custom_alu/mult/Q_reg[11]_i_1_n_2 ,\custom_alu/mult/Q_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[43] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[42] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[41] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[40] }),
        .O({\custom_alu/mult/Q_reg[11]_i_1_n_4 ,\custom_alu/mult/Q_reg[11]_i_1_n_5 ,\custom_alu/mult/Q_reg[11]_i_1_n_6 ,\custom_alu/mult/Q_reg[11]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[11]_i_2_n_0 ,\custom_alu/mult/Q[11]_i_3_n_0 ,\custom_alu/mult/Q[11]_i_4_n_0 ,\custom_alu/mult/Q[11]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[11]_i_8 
       (.CI(\custom_alu/mult/Q_reg[5]_i_4_n_0 ),
        .CO({\custom_alu/mult/Q_reg[11]_i_8_n_0 ,\custom_alu/mult/Q_reg[11]_i_8_n_1 ,\custom_alu/mult/Q_reg[11]_i_8_n_2 ,\custom_alu/mult/Q_reg[11]_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[71] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[70] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[69] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[68] }),
        .O(\custom_alu/MULT [38:35]),
        .S({\custom_alu/mult/Q[11]_i_12_n_0 ,\custom_alu/mult/Q[11]_i_13_n_0 ,\custom_alu/mult/Q[11]_i_14_n_0 ,\custom_alu/mult/Q[11]_i_15_n_0 }));
  CARRY4 \custom_alu/mult/Q_reg[15]_i_1 
       (.CI(\custom_alu/mult/Q_reg[11]_i_1_n_0 ),
        .CO({\custom_alu/mult/Q_reg[15]_i_1_n_0 ,\custom_alu/mult/Q_reg[15]_i_1_n_1 ,\custom_alu/mult/Q_reg[15]_i_1_n_2 ,\custom_alu/mult/Q_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[47] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[46] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[45] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[44] }),
        .O({\custom_alu/mult/Q_reg[15]_i_1_n_4 ,\custom_alu/mult/Q_reg[15]_i_1_n_5 ,\custom_alu/mult/Q_reg[15]_i_1_n_6 ,\custom_alu/mult/Q_reg[15]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[15]_i_2_n_0 ,\custom_alu/mult/Q[15]_i_3_n_0 ,\custom_alu/mult/Q[15]_i_4_n_0 ,\custom_alu/mult/Q[15]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[15]_i_5 
       (.CI(\custom_alu/mult/Q_reg[11]_i_8_n_0 ),
        .CO({\custom_alu/mult/Q_reg[15]_i_5_n_0 ,\custom_alu/mult/Q_reg[15]_i_5_n_1 ,\custom_alu/mult/Q_reg[15]_i_5_n_2 ,\custom_alu/mult/Q_reg[15]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[75] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[74] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[73] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[72] }),
        .O(\custom_alu/MULT [42:39]),
        .S({\custom_alu/mult/Q[15]_i_8_n_0 ,\custom_alu/mult/Q[15]_i_9_n_0 ,\custom_alu/mult/Q[15]_i_10_n_0 ,\custom_alu/mult/Q[15]_i_11_n_0 }));
  CARRY4 \custom_alu/mult/Q_reg[19]_i_1 
       (.CI(\custom_alu/mult/Q_reg[15]_i_1_n_0 ),
        .CO({\custom_alu/mult/Q_reg[19]_i_1_n_0 ,\custom_alu/mult/Q_reg[19]_i_1_n_1 ,\custom_alu/mult/Q_reg[19]_i_1_n_2 ,\custom_alu/mult/Q_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[51] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[50] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[49] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[48] }),
        .O({\custom_alu/mult/Q_reg[19]_i_1_n_4 ,\custom_alu/mult/Q_reg[19]_i_1_n_5 ,\custom_alu/mult/Q_reg[19]_i_1_n_6 ,\custom_alu/mult/Q_reg[19]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[19]_i_2_n_0 ,\custom_alu/mult/Q[19]_i_3_n_0 ,\custom_alu/mult/Q[19]_i_4_n_0 ,\custom_alu/mult/Q[19]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[19]_i_6 
       (.CI(\custom_alu/mult/Q_reg[15]_i_5_n_0 ),
        .CO({\custom_alu/mult/Q_reg[19]_i_6_n_0 ,\custom_alu/mult/Q_reg[19]_i_6_n_1 ,\custom_alu/mult/Q_reg[19]_i_6_n_2 ,\custom_alu/mult/Q_reg[19]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[79] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[78] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[77] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[76] }),
        .O(\custom_alu/MULT [46:43]),
        .S({\custom_alu/mult/Q[19]_i_8_n_0 ,\custom_alu/mult/Q[19]_i_9_n_0 ,\custom_alu/mult/Q[19]_i_10_n_0 ,\custom_alu/mult/Q[19]_i_11_n_0 }));
  CARRY4 \custom_alu/mult/Q_reg[23]_i_1 
       (.CI(\custom_alu/mult/Q_reg[19]_i_1_n_0 ),
        .CO({\custom_alu/mult/Q_reg[23]_i_1_n_0 ,\custom_alu/mult/Q_reg[23]_i_1_n_1 ,\custom_alu/mult/Q_reg[23]_i_1_n_2 ,\custom_alu/mult/Q_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[55] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[54] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[53] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[52] }),
        .O({\custom_alu/mult/Q_reg[23]_i_1_n_4 ,\custom_alu/mult/Q_reg[23]_i_1_n_5 ,\custom_alu/mult/Q_reg[23]_i_1_n_6 ,\custom_alu/mult/Q_reg[23]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[23]_i_2_n_0 ,\custom_alu/mult/Q[23]_i_3_n_0 ,\custom_alu/mult/Q[23]_i_4_n_0 ,\custom_alu/mult/Q[23]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[23]_i_4 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/Q_reg[23]_i_4_n_0 ,\custom_alu/mult/Q_reg[23]_i_4_n_1 ,\custom_alu/mult/Q_reg[23]_i_4_n_2 ,\custom_alu/mult/Q_reg[23]_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[51] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[50] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[49] ,\<const0> }),
        .O(\custom_alu/MULT [18:15]),
        .S({\custom_alu/mult/Q[23]_i_8_n_0 ,\custom_alu/mult/Q[23]_i_9_n_0 ,\custom_alu/mult/Q[23]_i_10_n_0 ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[48] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[23]_i_5 
       (.CI(\custom_alu/mult/Q_reg[19]_i_6_n_0 ),
        .CO({\custom_alu/mult/Q_reg[23]_i_5_n_0 ,\custom_alu/mult/Q_reg[23]_i_5_n_1 ,\custom_alu/mult/Q_reg[23]_i_5_n_2 ,\custom_alu/mult/Q_reg[23]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[81] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[80] }),
        .O(\custom_alu/MULT [50:47]),
        .S({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[83] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[82] ,\custom_alu/mult/Q[23]_i_11_n_0 ,\custom_alu/mult/Q[23]_i_12_n_0 }));
  CARRY4 \custom_alu/mult/Q_reg[27]_i_1 
       (.CI(\custom_alu/mult/Q_reg[23]_i_1_n_0 ),
        .CO({\custom_alu/mult/Q_reg[27]_i_1_n_0 ,\custom_alu/mult/Q_reg[27]_i_1_n_1 ,\custom_alu/mult/Q_reg[27]_i_1_n_2 ,\custom_alu/mult/Q_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[59] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[58] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[57] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[56] }),
        .O({\custom_alu/mult/Q_reg[27]_i_1_n_4 ,\custom_alu/mult/Q_reg[27]_i_1_n_5 ,\custom_alu/mult/Q_reg[27]_i_1_n_6 ,\custom_alu/mult/Q_reg[27]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[27]_i_2_n_0 ,\custom_alu/mult/Q[27]_i_3_n_0 ,\custom_alu/mult/Q[27]_i_4_n_0 ,\custom_alu/mult/Q[27]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[27]_i_4 
       (.CI(\custom_alu/mult/Q_reg[23]_i_4_n_0 ),
        .CO({\custom_alu/mult/Q_reg[27]_i_4_n_0 ,\custom_alu/mult/Q_reg[27]_i_4_n_1 ,\custom_alu/mult/Q_reg[27]_i_4_n_2 ,\custom_alu/mult/Q_reg[27]_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[55] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[54] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[53] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[52] }),
        .O(\custom_alu/MULT [22:19]),
        .S({\custom_alu/mult/Q[27]_i_9_n_0 ,\custom_alu/mult/Q[27]_i_10_n_0 ,\custom_alu/mult/Q[27]_i_11_n_0 ,\custom_alu/mult/Q[27]_i_12_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[27]_i_5 
       (.CI(\custom_alu/mult/Q_reg[23]_i_5_n_0 ),
        .CO({\custom_alu/mult/Q_reg[27]_i_5_n_0 ,\custom_alu/mult/Q_reg[27]_i_5_n_1 ,\custom_alu/mult/Q_reg[27]_i_5_n_2 ,\custom_alu/mult/Q_reg[27]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/MULT [54:51]),
        .S({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[87] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[86] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[85] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[84] }));
  CARRY4 \custom_alu/mult/Q_reg[31]_i_1 
       (.CI(\custom_alu/mult/Q_reg[27]_i_1_n_0 ),
        .CO({\custom_alu/mult/Q_reg[31]_i_1_n_0 ,\custom_alu/mult/Q_reg[31]_i_1_n_1 ,\custom_alu/mult/Q_reg[31]_i_1_n_2 ,\custom_alu/mult/Q_reg[31]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[63] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[62] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[61] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[60] }),
        .O({\custom_alu/mult/Q_reg[31]_i_1_n_4 ,\custom_alu/mult/Q_reg[31]_i_1_n_5 ,\custom_alu/mult/Q_reg[31]_i_1_n_6 ,\custom_alu/mult/Q_reg[31]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[31]_i_2_n_0 ,\custom_alu/mult/Q[31]_i_3_n_0 ,\custom_alu/mult/Q[31]_i_4_n_0 ,\custom_alu/mult/Q[31]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[31]_i_8 
       (.CI(\custom_alu/mult/Q_reg[27]_i_4_n_0 ),
        .CO({\custom_alu/mult/Q_reg[31]_i_8_n_0 ,\custom_alu/mult/Q_reg[31]_i_8_n_1 ,\custom_alu/mult/Q_reg[31]_i_8_n_2 ,\custom_alu/mult/Q_reg[31]_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[59] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[58] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[57] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[56] }),
        .O(\custom_alu/MULT [26:23]),
        .S({\custom_alu/mult/Q[31]_i_15_n_0 ,\custom_alu/mult/Q[31]_i_16_n_0 ,\custom_alu/mult/Q[31]_i_17_n_0 ,\custom_alu/mult/Q[31]_i_18_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[31]_i_9 
       (.CI(\custom_alu/mult/Q_reg[27]_i_5_n_0 ),
        .CO({\custom_alu/mult/Q_reg[31]_i_9_n_0 ,\custom_alu/mult/Q_reg[31]_i_9_n_1 ,\custom_alu/mult/Q_reg[31]_i_9_n_2 ,\custom_alu/mult/Q_reg[31]_i_9_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/MULT [58:55]),
        .S({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[91] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[90] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[89] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[88] }));
  CARRY4 \custom_alu/mult/Q_reg[32]_i_1 
       (.CI(\custom_alu/mult/Q_reg[31]_i_1_n_0 ),
        .CO(\custom_alu/mult/Q_reg[32]_i_1_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[35]_i_5 
       (.CI(\custom_alu/mult/Q_reg[31]_i_9_n_0 ),
        .CO({\custom_alu/mult/Q_reg[35]_i_5_n_0 ,\custom_alu/mult/Q_reg[35]_i_5_n_1 ,\custom_alu/mult/Q_reg[35]_i_5_n_2 ,\custom_alu/mult/Q_reg[35]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/MULT [62:59]),
        .S({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[95] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[94] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[93] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[92] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[35]_i_6 
       (.CI(\custom_alu/mult/Q_reg[31]_i_8_n_0 ),
        .CO({\custom_alu/mult/Q_reg[35]_i_6_n_0 ,\custom_alu/mult/Q_reg[35]_i_6_n_1 ,\custom_alu/mult/Q_reg[35]_i_6_n_2 ,\custom_alu/mult/Q_reg[35]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[63] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[62] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[61] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[60] }),
        .O(\custom_alu/MULT [30:27]),
        .S({\custom_alu/mult/Q[35]_i_12_n_0 ,\custom_alu/mult/Q[35]_i_13_n_0 ,\custom_alu/mult/Q[35]_i_14_n_0 ,\custom_alu/mult/Q[35]_i_15_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[36]_i_5 
       (.CI(\custom_alu/mult/Q_reg[35]_i_5_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/MULT [63]),
        .S({\<const0> ,\<const0> ,\<const0> ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[96] }));
  CARRY4 \custom_alu/mult/Q_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/Q_reg[3]_i_1_n_0 ,\custom_alu/mult/Q_reg[3]_i_1_n_1 ,\custom_alu/mult/Q_reg[3]_i_1_n_2 ,\custom_alu/mult/Q_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[35] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[34] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[33] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[32] }),
        .O({\custom_alu/mult/Q_reg[3]_i_1_n_4 ,\custom_alu/mult/Q_reg[3]_i_1_n_5 ,\custom_alu/mult/Q_reg[3]_i_1_n_6 ,\custom_alu/mult/Q_reg[3]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[3]_i_2_n_0 ,\custom_alu/mult/Q[3]_i_3_n_0 ,\custom_alu/mult/Q[3]_i_4_n_0 ,\custom_alu/mult/Q[3]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/Q_reg[5]_i_4 
       (.CI(\custom_alu/mult/Q_reg[35]_i_6_n_0 ),
        .CO({\custom_alu/mult/Q_reg[5]_i_4_n_0 ,\custom_alu/mult/Q_reg[5]_i_4_n_1 ,\custom_alu/mult/Q_reg[5]_i_4_n_2 ,\custom_alu/mult/Q_reg[5]_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[67] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[66] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[65] ,\custom_alu/mult/FF_MULT_1/Q_reg_n_0_[64] }),
        .O(\custom_alu/MULT [34:31]),
        .S({\custom_alu/mult/Q[5]_i_6_n_0 ,\custom_alu/mult/Q[5]_i_7_n_0 ,\custom_alu/mult/Q[5]_i_8_n_0 ,\custom_alu/mult/Q[5]_i_9_n_0 }));
  CARRY4 \custom_alu/mult/Q_reg[7]_i_1 
       (.CI(\custom_alu/mult/Q_reg[3]_i_1_n_0 ),
        .CO({\custom_alu/mult/Q_reg[7]_i_1_n_0 ,\custom_alu/mult/Q_reg[7]_i_1_n_1 ,\custom_alu/mult/Q_reg[7]_i_1_n_2 ,\custom_alu/mult/Q_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[39] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[38] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[37] ,\custom_alu/mult/FF_MULT_0/Q_reg_n_0_[36] }),
        .O({\custom_alu/mult/Q_reg[7]_i_1_n_4 ,\custom_alu/mult/Q_reg[7]_i_1_n_5 ,\custom_alu/mult/Q_reg[7]_i_1_n_6 ,\custom_alu/mult/Q_reg[7]_i_1_n_7 }),
        .S({\custom_alu/mult/Q[7]_i_2_n_0 ,\custom_alu/mult/Q[7]_i_3_n_0 ,\custom_alu/mult/Q[7]_i_4_n_0 ,\custom_alu/mult/Q[7]_i_5_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [0]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [10]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [11]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [12]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [13]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [14]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [15]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [0]),
        .Q(\custom_alu/mult/p_0_in [0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [1]),
        .Q(\custom_alu/mult/p_0_in [1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [2]),
        .Q(\custom_alu/mult/p_0_in [2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [3]),
        .Q(\custom_alu/mult/p_0_in [3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [1]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [4]),
        .Q(\custom_alu/mult/p_0_in [4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [5]),
        .Q(\custom_alu/mult/p_0_in [5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [6]),
        .Q(\custom_alu/mult/p_0_in [6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [7]),
        .Q(\custom_alu/mult/p_0_in [7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [8]),
        .Q(\custom_alu/mult/p_0_in [8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [9]),
        .Q(\custom_alu/mult/p_0_in [9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [10]),
        .Q(\custom_alu/mult/p_0_in [10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [11]),
        .Q(\custom_alu/mult/p_0_in [11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [12]),
        .Q(\custom_alu/mult/p_0_in [12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [13]),
        .Q(\custom_alu/mult/p_0_in [13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [2]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [14]),
        .Q(\custom_alu/mult/p_0_in [14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM2 [15]),
        .Q(\custom_alu/mult/p_0_in [15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [0]),
        .Q(\custom_alu/mult/p_1_in [0]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [1]),
        .Q(\custom_alu/mult/p_1_in [1]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [2]),
        .Q(\custom_alu/mult/p_1_in [2]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [3]),
        .Q(\custom_alu/mult/p_1_in [3]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [4]),
        .Q(\custom_alu/mult/p_1_in [4]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [5]),
        .Q(\custom_alu/mult/p_1_in [5]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [6]),
        .Q(\custom_alu/mult/p_1_in [6]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [7]),
        .Q(\custom_alu/mult/p_1_in [7]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [3]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [8]),
        .Q(\custom_alu/mult/p_1_in [8]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [9]),
        .Q(\custom_alu/mult/p_1_in [9]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [10]),
        .Q(\custom_alu/mult/p_1_in [10]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [11]),
        .Q(\custom_alu/mult/p_1_in [11]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [12]),
        .Q(\custom_alu/mult/p_1_in [12]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [13]),
        .Q(\custom_alu/mult/p_1_in [13]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [14]),
        .Q(\custom_alu/mult/p_1_in [14]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1 [15]),
        .Q(\custom_alu/mult/p_1_in [15]),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [4]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [7]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [8]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [9]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [10]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [11]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [5]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [12]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [13]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [14]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM0 [15]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[63] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [6]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [7]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [8]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_0/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM3 [9]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[9] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [0]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [10]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [11]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [12]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [13]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [14]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [15]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [16]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[16] ),
        .R(RST0));
  (* srl_bus_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/PSUM0 [0]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/PSUM0 [1]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/PSUM0 [2]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [1]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[1] ),
        .R(RST0));
  (* srl_bus_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/PSUM0 [3]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/PSUM0 [4]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/PSUM0 [5]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/PSUM0 [6]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[55] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[56] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[57] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[58] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[59] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[60] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [2]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[61] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[62] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[63] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[0] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[1] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[2] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[3] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[4] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[5] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[6] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [3]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[7] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[8] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[9] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[10] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[11] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[12] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[13] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[14] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_0/FF_MULT_0/Q_reg_n_0_[15] ),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [4]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [5]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [6]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [7]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [8]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_0/FF_MULT_1/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/PSUM1_2 [9]),
        .Q(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[9] ),
        .R(RST0));
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__0_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM0__0_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM0__0_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM0__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry_i_1__2_n_0,PSUM0__0_carry_i_2__0_n_0,PSUM0__0_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM0__0_carry_n_4 ,\custom_alu/mult/PSUM0 [2:0]}),
        .S({PSUM0__0_carry_i_4__0_n_0,PSUM0__0_carry_i_5__0_n_0,PSUM0__0_carry_i_6__2_n_0,PSUM0__0_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__0_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM0__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry__0_i_1__2_n_0,PSUM0__0_carry__0_i_2__2_n_0,PSUM0__0_carry__0_i_3__0_n_0,PSUM0__0_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_7 }),
        .S({PSUM0__0_carry__0_i_5__2_n_0,PSUM0__0_carry__0_i_6__2_n_0,PSUM0__0_carry__0_i_7__0_n_0,PSUM0__0_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__0_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM0__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__0_carry__1_i_1__2_n_0,PSUM0__0_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__0_carry__1_i_3__2_n_0,PSUM0__0_carry__1_i_4__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__30_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM0__30_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM0__30_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM0__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry_i_1__0_n_0,PSUM0__30_carry_i_2__2_n_0,PSUM0__30_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM0__30_carry_n_4 ,\custom_alu/mult/mult16_0/PSUM0__30_carry_n_5 ,\custom_alu/mult/mult16_0/PSUM0__30_carry_n_6 ,\custom_alu/mult/mult16_0/PSUM0__30_carry_n_7 }),
        .S({PSUM0__30_carry_i_4__0_n_0,PSUM0__30_carry_i_5__2_n_0,PSUM0__30_carry_i_6__2_n_0,PSUM0__30_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__30_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM0__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry__0_i_1__2_n_0,PSUM0__30_carry__0_i_2_n_0,PSUM0__30_carry__0_i_3__2_n_0,PSUM0__30_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_7 }),
        .S({PSUM0__30_carry__0_i_5__0_n_0,PSUM0__30_carry__0_i_6_n_0,PSUM0__30_carry__0_i_7_n_0,PSUM0__30_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__30_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM0__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM0__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__30_carry__1_i_1__2_n_0,PSUM0__30_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM0__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__30_carry__1_i_3__2_n_0,PSUM0__30_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__60_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM0__60_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM0__60_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM0__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry_i_1__2_n_0,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM0__0_carry__0_n_7 ,\custom_alu/mult/mult16_0/PSUM0__0_carry_n_4 }),
        .O(\custom_alu/mult/PSUM0 [6:3]),
        .S({PSUM0__60_carry_i_2__2_n_0,PSUM0__60_carry_i_3__2_n_0,PSUM0__60_carry_i_4__2_n_0,PSUM0__60_carry_i_5__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__60_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM0__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__0_i_1__2_n_0,PSUM0__60_carry__0_i_2__2_n_0,PSUM0__60_carry__0_i_3__2_n_0,PSUM0__60_carry__0_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM0 [10:7]),
        .S({PSUM0__60_carry__0_i_5__2_n_0,PSUM0__60_carry__0_i_6__2_n_0,PSUM0__60_carry__0_i_7__2_n_0,PSUM0__60_carry__0_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__60_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM0__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_0 ,\custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_1 ,\custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_2 ,\custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__1_i_1__2_n_0,PSUM0__60_carry__1_i_2__0_n_0,PSUM0__60_carry__1_i_3__2_n_0,PSUM0__60_carry__1_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM0 [14:11]),
        .S({PSUM0__60_carry__1_i_5__0_n_0,PSUM0__60_carry__1_i_6__0_n_0,PSUM0__60_carry__1_i_7__0_n_0,PSUM0__60_carry__1_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM0__60_carry__2 
       (.CI(\custom_alu/mult/mult16_0/PSUM0__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/PSUM0 [15]),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM0__60_carry__2_i_1__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__0_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM1__0_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM1__0_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM1__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry_i_1__2_n_0,PSUM1__0_carry_i_2__2_n_0,PSUM1__0_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM1__0_carry_n_4 ,\custom_alu/mult/PSUM1 [2:0]}),
        .S({PSUM1__0_carry_i_4__2_n_0,PSUM1__0_carry_i_5__2_n_0,PSUM1__0_carry_i_6__2_n_0,PSUM1__0_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__0_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM1__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry__0_i_1__2_n_0,PSUM1__0_carry__0_i_2__2_n_0,PSUM1__0_carry__0_i_3__2_n_0,PSUM1__0_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_7 }),
        .S({PSUM1__0_carry__0_i_5__2_n_0,PSUM1__0_carry__0_i_6__2_n_0,PSUM1__0_carry__0_i_7__2_n_0,PSUM1__0_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__0_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM1__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__0_carry__1_i_1__2_n_0,PSUM1__0_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__0_carry__1_i_3__2_n_0,PSUM1__0_carry__1_i_4__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__30_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM1__30_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM1__30_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM1__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry_i_1__2_n_0,PSUM1__30_carry_i_2__2_n_0,PSUM1__30_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM1__30_carry_n_4 ,\custom_alu/mult/mult16_0/PSUM1__30_carry_n_5 ,\custom_alu/mult/mult16_0/PSUM1__30_carry_n_6 ,\custom_alu/mult/mult16_0/PSUM1__30_carry_n_7 }),
        .S({PSUM1__30_carry_i_4__2_n_0,PSUM1__30_carry_i_5__2_n_0,PSUM1__30_carry_i_6__2_n_0,PSUM1__30_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__30_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM1__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry__0_i_1__2_n_0,PSUM1__30_carry__0_i_2__2_n_0,PSUM1__30_carry__0_i_3__2_n_0,PSUM1__30_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_7 }),
        .S({PSUM1__30_carry__0_i_5__2_n_0,PSUM1__30_carry__0_i_6__2_n_0,PSUM1__30_carry__0_i_7__2_n_0,PSUM1__30_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__30_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM1__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM1__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__30_carry__1_i_1__2_n_0,PSUM1__30_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM1__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__30_carry__1_i_3__2_n_0,PSUM1__30_carry__1_i_4__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__60_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM1__60_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM1__60_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM1__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry_i_1__2_n_0,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM1__0_carry__0_n_7 ,\custom_alu/mult/mult16_0/PSUM1__0_carry_n_4 }),
        .O(\custom_alu/mult/PSUM1 [6:3]),
        .S({PSUM1__60_carry_i_2__2_n_0,PSUM1__60_carry_i_3__2_n_0,PSUM1__60_carry_i_4__2_n_0,PSUM1__60_carry_i_5__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__60_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM1__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__0_i_1__2_n_0,PSUM1__60_carry__0_i_2__2_n_0,PSUM1__60_carry__0_i_3__2_n_0,PSUM1__60_carry__0_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM1 [10:7]),
        .S({PSUM1__60_carry__0_i_5__2_n_0,PSUM1__60_carry__0_i_6__2_n_0,PSUM1__60_carry__0_i_7__2_n_0,PSUM1__60_carry__0_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__60_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM1__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_0 ,\custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_1 ,\custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_2 ,\custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__1_i_1__2_n_0,PSUM1__60_carry__1_i_2__2_n_0,PSUM1__60_carry__1_i_3__2_n_0,PSUM1__60_carry__1_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM1 [14:11]),
        .S({PSUM1__60_carry__1_i_5__2_n_0,PSUM1__60_carry__1_i_6__2_n_0,PSUM1__60_carry__1_i_7__2_n_0,PSUM1__60_carry__1_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM1__60_carry__2 
       (.CI(\custom_alu/mult/mult16_0/PSUM1__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/PSUM1 [15]),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM1__60_carry__2_i_1__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__0_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM2__0_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM2__0_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM2__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry_i_1__2_n_0,PSUM2__0_carry_i_2__2_n_0,PSUM2__0_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM2__0_carry_n_4 ,\custom_alu/mult/PSUM2 [2:0]}),
        .S({PSUM2__0_carry_i_4__2_n_0,PSUM2__0_carry_i_5__2_n_0,PSUM2__0_carry_i_6__2_n_0,PSUM2__0_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__0_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM2__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry__0_i_1__2_n_0,PSUM2__0_carry__0_i_2__2_n_0,PSUM2__0_carry__0_i_3__2_n_0,PSUM2__0_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_7 }),
        .S({PSUM2__0_carry__0_i_5__2_n_0,PSUM2__0_carry__0_i_6__2_n_0,PSUM2__0_carry__0_i_7__2_n_0,PSUM2__0_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__0_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM2__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__0_carry__1_i_1__2_n_0,PSUM2__0_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__0_carry__1_i_3__2_n_0,PSUM2__0_carry__1_i_4__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__30_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM2__30_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM2__30_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM2__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry_i_1__2_n_0,PSUM2__30_carry_i_2__2_n_0,PSUM2__30_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM2__30_carry_n_4 ,\custom_alu/mult/mult16_0/PSUM2__30_carry_n_5 ,\custom_alu/mult/mult16_0/PSUM2__30_carry_n_6 ,\custom_alu/mult/mult16_0/PSUM2__30_carry_n_7 }),
        .S({PSUM2__30_carry_i_4__2_n_0,PSUM2__30_carry_i_5__2_n_0,PSUM2__30_carry_i_6__2_n_0,PSUM2__30_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__30_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM2__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry__0_i_1__2_n_0,PSUM2__30_carry__0_i_2__2_n_0,PSUM2__30_carry__0_i_3__2_n_0,PSUM2__30_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_7 }),
        .S({PSUM2__30_carry__0_i_5__2_n_0,PSUM2__30_carry__0_i_6__2_n_0,PSUM2__30_carry__0_i_7__2_n_0,PSUM2__30_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__30_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM2__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM2__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__30_carry__1_i_1__2_n_0,PSUM2__30_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM2__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__30_carry__1_i_3__2_n_0,PSUM2__30_carry__1_i_4__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__60_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM2__60_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM2__60_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM2__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry_i_1__2_n_0,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM2__0_carry__0_n_7 ,\custom_alu/mult/mult16_0/PSUM2__0_carry_n_4 }),
        .O(\custom_alu/mult/PSUM2 [6:3]),
        .S({PSUM2__60_carry_i_2__2_n_0,PSUM2__60_carry_i_3__2_n_0,PSUM2__60_carry_i_4__2_n_0,PSUM2__60_carry_i_5__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__60_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM2__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__0_i_1__2_n_0,PSUM2__60_carry__0_i_2__2_n_0,PSUM2__60_carry__0_i_3__2_n_0,PSUM2__60_carry__0_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM2 [10:7]),
        .S({PSUM2__60_carry__0_i_5__2_n_0,PSUM2__60_carry__0_i_6__2_n_0,PSUM2__60_carry__0_i_7__2_n_0,PSUM2__60_carry__0_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__60_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM2__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_0 ,\custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_1 ,\custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_2 ,\custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__1_i_1__2_n_0,PSUM2__60_carry__1_i_2__2_n_0,PSUM2__60_carry__1_i_3__2_n_0,PSUM2__60_carry__1_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM2 [14:11]),
        .S({PSUM2__60_carry__1_i_5__2_n_0,PSUM2__60_carry__1_i_6__2_n_0,PSUM2__60_carry__1_i_7__2_n_0,PSUM2__60_carry__1_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM2__60_carry__2 
       (.CI(\custom_alu/mult/mult16_0/PSUM2__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/PSUM2 [15]),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM2__60_carry__2_i_1__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__0_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM3__0_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM3__0_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM3__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry_i_1__2_n_0,PSUM3__0_carry_i_2__0_n_0,PSUM3__0_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM3__0_carry_n_4 ,\custom_alu/mult/PSUM3 [2:0]}),
        .S({PSUM3__0_carry_i_4__0_n_0,PSUM3__0_carry_i_5__0_n_0,PSUM3__0_carry_i_6__2_n_0,PSUM3__0_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__0_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM3__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry__0_i_1__2_n_0,PSUM3__0_carry__0_i_2__2_n_0,PSUM3__0_carry__0_i_3__0_n_0,PSUM3__0_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_7 }),
        .S({PSUM3__0_carry__0_i_5__2_n_0,PSUM3__0_carry__0_i_6__2_n_0,PSUM3__0_carry__0_i_7__0_n_0,PSUM3__0_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__0_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM3__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__0_carry__1_i_1__2_n_0,PSUM3__0_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__0_carry__1_i_3__2_n_0,PSUM3__0_carry__1_i_4__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__30_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM3__30_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM3__30_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM3__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry_i_1__0_n_0,PSUM3__30_carry_i_2__2_n_0,PSUM3__30_carry_i_3__2_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_0/PSUM3__30_carry_n_4 ,\custom_alu/mult/mult16_0/PSUM3__30_carry_n_5 ,\custom_alu/mult/mult16_0/PSUM3__30_carry_n_6 ,\custom_alu/mult/mult16_0/PSUM3__30_carry_n_7 }),
        .S({PSUM3__30_carry_i_4__0_n_0,PSUM3__30_carry_i_5__2_n_0,PSUM3__30_carry_i_6__2_n_0,PSUM3__30_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__30_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM3__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry__0_i_1__2_n_0,PSUM3__30_carry__0_i_2__0_n_0,PSUM3__30_carry__0_i_3__2_n_0,PSUM3__30_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_4 ,\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_5 ,\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_7 }),
        .S({PSUM3__30_carry__0_i_5__0_n_0,PSUM3__30_carry__0_i_6__0_n_0,PSUM3__30_carry__0_i_7__0_n_0,PSUM3__30_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__30_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM3__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_0/PSUM3__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__30_carry__1_i_1__2_n_0,PSUM3__30_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_6 ,\custom_alu/mult/mult16_0/PSUM3__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__30_carry__1_i_3__2_n_0,PSUM3__30_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__60_carry_n_0 ,\custom_alu/mult/mult16_0/PSUM3__60_carry_n_1 ,\custom_alu/mult/mult16_0/PSUM3__60_carry_n_2 ,\custom_alu/mult/mult16_0/PSUM3__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry_i_1__2_n_0,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_0/PSUM3__0_carry__0_n_7 ,\custom_alu/mult/mult16_0/PSUM3__0_carry_n_4 }),
        .O(\custom_alu/mult/PSUM3 [6:3]),
        .S({PSUM3__60_carry_i_2__2_n_0,PSUM3__60_carry_i_3__2_n_0,PSUM3__60_carry_i_4__2_n_0,PSUM3__60_carry_i_5__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__60_carry__0 
       (.CI(\custom_alu/mult/mult16_0/PSUM3__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_0 ,\custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_1 ,\custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_2 ,\custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__0_i_1__2_n_0,PSUM3__60_carry__0_i_2__2_n_0,PSUM3__60_carry__0_i_3__2_n_0,PSUM3__60_carry__0_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM3 [10:7]),
        .S({PSUM3__60_carry__0_i_5__2_n_0,PSUM3__60_carry__0_i_6__2_n_0,PSUM3__60_carry__0_i_7__2_n_0,PSUM3__60_carry__0_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__60_carry__1 
       (.CI(\custom_alu/mult/mult16_0/PSUM3__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_0 ,\custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_1 ,\custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_2 ,\custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__1_i_1__2_n_0,PSUM3__60_carry__1_i_2__0_n_0,PSUM3__60_carry__1_i_3__2_n_0,PSUM3__60_carry__1_i_4__2_n_0}),
        .O(\custom_alu/mult/PSUM3 [14:11]),
        .S({PSUM3__60_carry__1_i_5__0_n_0,PSUM3__60_carry__1_i_6__0_n_0,PSUM3__60_carry__1_i_7__0_n_0,PSUM3__60_carry__1_i_8__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/PSUM3__60_carry__2 
       (.CI(\custom_alu/mult/mult16_0/PSUM3__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/PSUM3 [15]),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM3__60_carry__2_i_1__0_n_0}));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[106]_i_2 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[27] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[2] ),
        .O(\custom_alu/mult/mult16_0/Q[106]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[106]_i_3 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[26] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[1] ),
        .O(\custom_alu/mult/mult16_0/Q[106]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[106]_i_4 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[25] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[0] ),
        .O(\custom_alu/mult/mult16_0/Q[106]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[110]_i_2 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[31] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[6] ),
        .O(\custom_alu/mult/mult16_0/Q[110]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[110]_i_3 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[30] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[5] ),
        .O(\custom_alu/mult/mult16_0/Q[110]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[110]_i_4 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[29] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[4] ),
        .O(\custom_alu/mult/mult16_0/Q[110]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[110]_i_5 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[28] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[3] ),
        .O(\custom_alu/mult/mult16_0/Q[110]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[114]_i_2 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[10] ),
        .O(\custom_alu/mult/mult16_0/Q[114]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[114]_i_3 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[9] ),
        .O(\custom_alu/mult/mult16_0/Q[114]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[114]_i_4 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[8] ),
        .O(\custom_alu/mult/mult16_0/Q[114]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[114]_i_5 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[7] ),
        .O(\custom_alu/mult/mult16_0/Q[114]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[118]_i_2 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[14] ),
        .O(\custom_alu/mult/mult16_0/Q[118]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[118]_i_3 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[13] ),
        .O(\custom_alu/mult/mult16_0/Q[118]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[118]_i_4 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[12] ),
        .O(\custom_alu/mult/mult16_0/Q[118]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[118]_i_5 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[11] ),
        .O(\custom_alu/mult/mult16_0/Q[118]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[11]_i_2 
       (.I0(\custom_alu/mult/p_1_in [11]),
        .I1(\custom_alu/mult/p_0_in [11]),
        .O(\custom_alu/mult/mult16_0/Q[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[11]_i_3 
       (.I0(\custom_alu/mult/p_1_in [10]),
        .I1(\custom_alu/mult/p_0_in [10]),
        .O(\custom_alu/mult/mult16_0/Q[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[11]_i_4 
       (.I0(\custom_alu/mult/p_1_in [9]),
        .I1(\custom_alu/mult/p_0_in [9]),
        .O(\custom_alu/mult/mult16_0/Q[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[11]_i_5 
       (.I0(\custom_alu/mult/p_1_in [8]),
        .I1(\custom_alu/mult/p_0_in [8]),
        .O(\custom_alu/mult/mult16_0/Q[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[122]_i_2 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/mult16_0/Q[122]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[122]_i_3 
       (.I0(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[15] ),
        .O(\custom_alu/mult/mult16_0/Q[122]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[15]_i_2 
       (.I0(\custom_alu/mult/p_1_in [15]),
        .I1(\custom_alu/mult/p_0_in [15]),
        .O(\custom_alu/mult/mult16_0/Q[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[15]_i_3 
       (.I0(\custom_alu/mult/p_1_in [14]),
        .I1(\custom_alu/mult/p_0_in [14]),
        .O(\custom_alu/mult/mult16_0/Q[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[15]_i_4 
       (.I0(\custom_alu/mult/p_1_in [13]),
        .I1(\custom_alu/mult/p_0_in [13]),
        .O(\custom_alu/mult/mult16_0/Q[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[15]_i_5 
       (.I0(\custom_alu/mult/p_1_in [12]),
        .I1(\custom_alu/mult/p_0_in [12]),
        .O(\custom_alu/mult/mult16_0/Q[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[3]_i_2 
       (.I0(\custom_alu/mult/p_1_in [3]),
        .I1(\custom_alu/mult/p_0_in [3]),
        .O(\custom_alu/mult/mult16_0/Q[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[3]_i_3 
       (.I0(\custom_alu/mult/p_1_in [2]),
        .I1(\custom_alu/mult/p_0_in [2]),
        .O(\custom_alu/mult/mult16_0/Q[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[3]_i_4 
       (.I0(\custom_alu/mult/p_1_in [1]),
        .I1(\custom_alu/mult/p_0_in [1]),
        .O(\custom_alu/mult/mult16_0/Q[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[3]_i_5 
       (.I0(\custom_alu/mult/p_1_in [0]),
        .I1(\custom_alu/mult/p_0_in [0]),
        .O(\custom_alu/mult/mult16_0/Q[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[7]_i_2 
       (.I0(\custom_alu/mult/p_1_in [7]),
        .I1(\custom_alu/mult/p_0_in [7]),
        .O(\custom_alu/mult/mult16_0/Q[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[7]_i_3 
       (.I0(\custom_alu/mult/p_1_in [6]),
        .I1(\custom_alu/mult/p_0_in [6]),
        .O(\custom_alu/mult/mult16_0/Q[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[7]_i_4 
       (.I0(\custom_alu/mult/p_1_in [5]),
        .I1(\custom_alu/mult/p_0_in [5]),
        .O(\custom_alu/mult/mult16_0/Q[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_0/Q[7]_i_5 
       (.I0(\custom_alu/mult/p_1_in [4]),
        .I1(\custom_alu/mult/p_0_in [4]),
        .O(\custom_alu/mult/mult16_0/Q[7]_i_5_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[106]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[27] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[26] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[25] ,\<const0> }),
        .O(\custom_alu/mult/PSUM0_1_2_3 [10:7]),
        .S({\custom_alu/mult/mult16_0/Q[106]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[106]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[106]_i_4_n_0 ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[24] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[110]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[106]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[31] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[30] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[29] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[28] }),
        .O(\custom_alu/mult/PSUM0_1_2_3 [14:11]),
        .S({\custom_alu/mult/mult16_0/Q[110]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[110]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[110]_i_4_n_0 ,\custom_alu/mult/mult16_0/Q[110]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[114]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[110]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[35] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[34] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[33] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[32] }),
        .O(\custom_alu/mult/PSUM0_1_2_3 [18:15]),
        .S({\custom_alu/mult/mult16_0/Q[114]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[114]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[114]_i_4_n_0 ,\custom_alu/mult/mult16_0/Q[114]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[118]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[114]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[39] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[38] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[37] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[36] }),
        .O(\custom_alu/mult/PSUM0_1_2_3 [22:19]),
        .S({\custom_alu/mult/mult16_0/Q[118]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[118]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[118]_i_4_n_0 ,\custom_alu/mult/mult16_0/Q[118]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[11]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/mult/p_1_in [11:8]),
        .O(\custom_alu/mult/PSUM1_2 [11:8]),
        .S({\custom_alu/mult/mult16_0/Q[11]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[11]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[11]_i_4_n_0 ,\custom_alu/mult/mult16_0/Q[11]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[122]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[118]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[41] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[40] }),
        .O(\custom_alu/mult/PSUM0_1_2_3 [26:23]),
        .S({\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[43] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[42] ,\custom_alu/mult/mult16_0/Q[122]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[122]_i_3_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[126]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[122]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/PSUM0_1_2_3 [30:27]),
        .S({\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[47] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[46] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[45] ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[44] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[127]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[126]_i_1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/PSUM0_1_2_3 [31]),
        .S({\<const0> ,\<const0> ,\<const0> ,\custom_alu/mult/mult16_0/FF_MULT_1/Q_reg_n_0_[48] }));
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[15]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[11]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/mult/p_1_in [15:12]),
        .O(\custom_alu/mult/PSUM1_2 [15:12]),
        .S({\custom_alu/mult/mult16_0/Q[15]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[15]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[15]_i_4_n_0 ,\custom_alu/mult/mult16_0/Q[15]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[16]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[15]_i_1_n_0 ),
        .CO(\custom_alu/mult/PSUM1_2 [16]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/mult/p_1_in [3:0]),
        .O(\custom_alu/mult/PSUM1_2 [3:0]),
        .S({\custom_alu/mult/mult16_0/Q[3]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[3]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[3]_i_4_n_0 ,\custom_alu/mult/mult16_0/Q[3]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_0/Q_reg[7]_i_1 
       (.CI(\custom_alu/mult/mult16_0/Q_reg[3]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_0 ,\custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_1 ,\custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_2 ,\custom_alu/mult/mult16_0/Q_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\custom_alu/mult/p_1_in [7:4]),
        .O(\custom_alu/mult/PSUM1_2 [7:4]),
        .S({\custom_alu/mult/mult16_0/Q[7]_i_2_n_0 ,\custom_alu/mult/mult16_0/Q[7]_i_3_n_0 ,\custom_alu/mult/mult16_0/Q[7]_i_4_n_0 ,\custom_alu/mult/mult16_0/Q[7]_i_5_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM2__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM1__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[49] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[49] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[50] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[50] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[51] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[51] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[52] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[52] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[53] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[53] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[54] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[54] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM0__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[63] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_0/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[9] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[16]_i_1_n_3 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[48] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[49] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[50] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[51] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[52] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[53] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[54] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[55] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[56] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[57] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[58] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[59] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[60] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[61] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[62] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[63] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[0] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[1] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[2] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[3] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[4] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[5] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[6] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[7] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[8] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[9] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[10] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[11] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[12] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[13] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[14] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[15] ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_1/FF_MULT_1/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[9] ),
        .R(RST0));
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__0_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM0__0_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM0__0_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM0__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry_i_1__1_n_0,PSUM0__0_carry_i_2__2_n_0,PSUM0__0_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM0__0_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM0__0_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM0__0_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM0__0_carry_n_7 }),
        .S({PSUM0__0_carry_i_4__2_n_0,PSUM0__0_carry_i_5__2_n_0,PSUM0__0_carry_i_6__1_n_0,PSUM0__0_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__0_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM0__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry__0_i_1__1_n_0,PSUM0__0_carry__0_i_2__1_n_0,PSUM0__0_carry__0_i_3__2_n_0,PSUM0__0_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_7 }),
        .S({PSUM0__0_carry__0_i_5__1_n_0,PSUM0__0_carry__0_i_6__1_n_0,PSUM0__0_carry__0_i_7__2_n_0,PSUM0__0_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__0_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM0__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__0_carry__1_i_1__1_n_0,PSUM0__0_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__0_carry__1_i_3__1_n_0,PSUM0__0_carry__1_i_4__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__30_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM0__30_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM0__30_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM0__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry_i_1__2_n_0,PSUM0__30_carry_i_2__1_n_0,PSUM0__30_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM0__30_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM0__30_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM0__30_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM0__30_carry_n_7 }),
        .S({PSUM0__30_carry_i_4__2_n_0,PSUM0__30_carry_i_5__1_n_0,PSUM0__30_carry_i_6__1_n_0,PSUM0__30_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__30_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM0__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry__0_i_1__1_n_0,PSUM0__30_carry__0_i_2__2_n_0,PSUM0__30_carry__0_i_3__1_n_0,PSUM0__30_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_7 }),
        .S({PSUM0__30_carry__0_i_5__2_n_0,PSUM0__30_carry__0_i_6__2_n_0,PSUM0__30_carry__0_i_7__2_n_0,PSUM0__30_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__30_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM0__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM0__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__30_carry__1_i_1__1_n_0,PSUM0__30_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM0__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__30_carry__1_i_3__1_n_0,PSUM0__30_carry__1_i_4__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__60_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM0__60_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM0__60_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM0__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry_i_1__1_n_0,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM0__0_carry__0_n_7 ,\custom_alu/mult/mult16_1/PSUM0__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_1/PSUM0__60_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM0__60_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM0__60_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM0__60_carry_n_7 }),
        .S({PSUM0__60_carry_i_2__1_n_0,PSUM0__60_carry_i_3__1_n_0,PSUM0__60_carry_i_4__1_n_0,PSUM0__60_carry_i_5__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__60_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM0__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__0_i_1__1_n_0,PSUM0__60_carry__0_i_2__1_n_0,PSUM0__60_carry__0_i_3__1_n_0,PSUM0__60_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_7 }),
        .S({PSUM0__60_carry__0_i_5__1_n_0,PSUM0__60_carry__0_i_6__1_n_0,PSUM0__60_carry__0_i_7__1_n_0,PSUM0__60_carry__0_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__60_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM0__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_0 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_1 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_2 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__1_i_1__1_n_0,PSUM0__60_carry__1_i_2__2_n_0,PSUM0__60_carry__1_i_3__1_n_0,PSUM0__60_carry__1_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_4 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_5 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_7 }),
        .S({PSUM0__60_carry__1_i_5__2_n_0,PSUM0__60_carry__1_i_6__2_n_0,PSUM0__60_carry__1_i_7__2_n_0,PSUM0__60_carry__1_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM0__60_carry__2 
       (.CI(\custom_alu/mult/mult16_1/PSUM0__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_1/PSUM0__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM0__60_carry__2_i_1__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__0_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM1__0_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM1__0_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM1__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry_i_1__1_n_0,PSUM1__0_carry_i_2__1_n_0,PSUM1__0_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM1__0_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM1__0_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM1__0_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM1__0_carry_n_7 }),
        .S({PSUM1__0_carry_i_4__1_n_0,PSUM1__0_carry_i_5__1_n_0,PSUM1__0_carry_i_6__1_n_0,PSUM1__0_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__0_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM1__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry__0_i_1__1_n_0,PSUM1__0_carry__0_i_2__1_n_0,PSUM1__0_carry__0_i_3__1_n_0,PSUM1__0_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_7 }),
        .S({PSUM1__0_carry__0_i_5__1_n_0,PSUM1__0_carry__0_i_6__1_n_0,PSUM1__0_carry__0_i_7__1_n_0,PSUM1__0_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__0_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM1__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__0_carry__1_i_1__1_n_0,PSUM1__0_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__0_carry__1_i_3__1_n_0,PSUM1__0_carry__1_i_4__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__30_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM1__30_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM1__30_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM1__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry_i_1__1_n_0,PSUM1__30_carry_i_2__1_n_0,PSUM1__30_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM1__30_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM1__30_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM1__30_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM1__30_carry_n_7 }),
        .S({PSUM1__30_carry_i_4__1_n_0,PSUM1__30_carry_i_5__1_n_0,PSUM1__30_carry_i_6__1_n_0,PSUM1__30_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__30_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM1__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry__0_i_1__1_n_0,PSUM1__30_carry__0_i_2__1_n_0,PSUM1__30_carry__0_i_3__1_n_0,PSUM1__30_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_7 }),
        .S({PSUM1__30_carry__0_i_5__1_n_0,PSUM1__30_carry__0_i_6__1_n_0,PSUM1__30_carry__0_i_7__1_n_0,PSUM1__30_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__30_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM1__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM1__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__30_carry__1_i_1__1_n_0,PSUM1__30_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM1__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__30_carry__1_i_3__1_n_0,PSUM1__30_carry__1_i_4__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__60_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM1__60_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM1__60_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM1__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry_i_1__1_n_0,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM1__0_carry__0_n_7 ,\custom_alu/mult/mult16_1/PSUM1__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_1/PSUM1__60_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM1__60_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM1__60_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM1__60_carry_n_7 }),
        .S({PSUM1__60_carry_i_2__1_n_0,PSUM1__60_carry_i_3__1_n_0,PSUM1__60_carry_i_4__1_n_0,PSUM1__60_carry_i_5__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__60_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM1__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__0_i_1__1_n_0,PSUM1__60_carry__0_i_2__1_n_0,PSUM1__60_carry__0_i_3__1_n_0,PSUM1__60_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_7 }),
        .S({PSUM1__60_carry__0_i_5__1_n_0,PSUM1__60_carry__0_i_6__1_n_0,PSUM1__60_carry__0_i_7__1_n_0,PSUM1__60_carry__0_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__60_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM1__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_0 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_1 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_2 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__1_i_1__1_n_0,PSUM1__60_carry__1_i_2__1_n_0,PSUM1__60_carry__1_i_3__1_n_0,PSUM1__60_carry__1_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_4 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_5 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_7 }),
        .S({PSUM1__60_carry__1_i_5__1_n_0,PSUM1__60_carry__1_i_6__1_n_0,PSUM1__60_carry__1_i_7__1_n_0,PSUM1__60_carry__1_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM1__60_carry__2 
       (.CI(\custom_alu/mult/mult16_1/PSUM1__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_1/PSUM1__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM1__60_carry__2_i_1__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__0_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM2__0_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM2__0_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM2__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry_i_1__1_n_0,PSUM2__0_carry_i_2__1_n_0,PSUM2__0_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM2__0_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM2__0_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM2__0_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM2__0_carry_n_7 }),
        .S({PSUM2__0_carry_i_4__1_n_0,PSUM2__0_carry_i_5__1_n_0,PSUM2__0_carry_i_6__1_n_0,PSUM2__0_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__0_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM2__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry__0_i_1__1_n_0,PSUM2__0_carry__0_i_2__1_n_0,PSUM2__0_carry__0_i_3__1_n_0,PSUM2__0_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_7 }),
        .S({PSUM2__0_carry__0_i_5__1_n_0,PSUM2__0_carry__0_i_6__1_n_0,PSUM2__0_carry__0_i_7__1_n_0,PSUM2__0_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__0_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM2__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__0_carry__1_i_1__1_n_0,PSUM2__0_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__0_carry__1_i_3__1_n_0,PSUM2__0_carry__1_i_4__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__30_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM2__30_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM2__30_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM2__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry_i_1__1_n_0,PSUM2__30_carry_i_2__1_n_0,PSUM2__30_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM2__30_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM2__30_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM2__30_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM2__30_carry_n_7 }),
        .S({PSUM2__30_carry_i_4__1_n_0,PSUM2__30_carry_i_5__1_n_0,PSUM2__30_carry_i_6__1_n_0,PSUM2__30_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__30_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM2__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry__0_i_1__1_n_0,PSUM2__30_carry__0_i_2__1_n_0,PSUM2__30_carry__0_i_3__1_n_0,PSUM2__30_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_7 }),
        .S({PSUM2__30_carry__0_i_5__1_n_0,PSUM2__30_carry__0_i_6__1_n_0,PSUM2__30_carry__0_i_7__1_n_0,PSUM2__30_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__30_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM2__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM2__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__30_carry__1_i_1__1_n_0,PSUM2__30_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM2__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__30_carry__1_i_3__1_n_0,PSUM2__30_carry__1_i_4__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__60_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM2__60_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM2__60_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM2__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry_i_1__1_n_0,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM2__0_carry__0_n_7 ,\custom_alu/mult/mult16_1/PSUM2__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_1/PSUM2__60_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM2__60_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM2__60_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM2__60_carry_n_7 }),
        .S({PSUM2__60_carry_i_2__1_n_0,PSUM2__60_carry_i_3__1_n_0,PSUM2__60_carry_i_4__1_n_0,PSUM2__60_carry_i_5__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__60_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM2__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__0_i_1__1_n_0,PSUM2__60_carry__0_i_2__1_n_0,PSUM2__60_carry__0_i_3__1_n_0,PSUM2__60_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_7 }),
        .S({PSUM2__60_carry__0_i_5__1_n_0,PSUM2__60_carry__0_i_6__1_n_0,PSUM2__60_carry__0_i_7__1_n_0,PSUM2__60_carry__0_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__60_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM2__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_0 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_1 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_2 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__1_i_1__1_n_0,PSUM2__60_carry__1_i_2__1_n_0,PSUM2__60_carry__1_i_3__1_n_0,PSUM2__60_carry__1_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_4 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_5 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_7 }),
        .S({PSUM2__60_carry__1_i_5__1_n_0,PSUM2__60_carry__1_i_6__1_n_0,PSUM2__60_carry__1_i_7__1_n_0,PSUM2__60_carry__1_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM2__60_carry__2 
       (.CI(\custom_alu/mult/mult16_1/PSUM2__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_1/PSUM2__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM2__60_carry__2_i_1__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__0_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM3__0_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM3__0_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM3__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry_i_1__1_n_0,PSUM3__0_carry_i_2__2_n_0,PSUM3__0_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM3__0_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM3__0_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM3__0_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM3__0_carry_n_7 }),
        .S({PSUM3__0_carry_i_4__2_n_0,PSUM3__0_carry_i_5__2_n_0,PSUM3__0_carry_i_6__1_n_0,PSUM3__0_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__0_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM3__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry__0_i_1__1_n_0,PSUM3__0_carry__0_i_2__1_n_0,PSUM3__0_carry__0_i_3__2_n_0,PSUM3__0_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_7 }),
        .S({PSUM3__0_carry__0_i_5__1_n_0,PSUM3__0_carry__0_i_6__1_n_0,PSUM3__0_carry__0_i_7__2_n_0,PSUM3__0_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__0_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM3__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__0_carry__1_i_1__1_n_0,PSUM3__0_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__0_carry__1_i_3__1_n_0,PSUM3__0_carry__1_i_4__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__30_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM3__30_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM3__30_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM3__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry_i_1__2_n_0,PSUM3__30_carry_i_2__1_n_0,PSUM3__30_carry_i_3__1_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_1/PSUM3__30_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM3__30_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM3__30_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM3__30_carry_n_7 }),
        .S({PSUM3__30_carry_i_4__2_n_0,PSUM3__30_carry_i_5__1_n_0,PSUM3__30_carry_i_6__1_n_0,PSUM3__30_carry_i_7_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__30_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM3__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry__0_i_1__1_n_0,PSUM3__30_carry__0_i_2__2_n_0,PSUM3__30_carry__0_i_3__1_n_0,PSUM3__30_carry__0_i_4__2_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_7 }),
        .S({PSUM3__30_carry__0_i_5__2_n_0,PSUM3__30_carry__0_i_6__2_n_0,PSUM3__30_carry__0_i_7__2_n_0,PSUM3__30_carry__0_i_8__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__30_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM3__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_1/PSUM3__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__30_carry__1_i_1__1_n_0,PSUM3__30_carry__1_i_2__2_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM3__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__30_carry__1_i_3__1_n_0,PSUM3__30_carry__1_i_4__2_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__60_carry_n_0 ,\custom_alu/mult/mult16_1/PSUM3__60_carry_n_1 ,\custom_alu/mult/mult16_1/PSUM3__60_carry_n_2 ,\custom_alu/mult/mult16_1/PSUM3__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry_i_1__1_n_0,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM3__0_carry__0_n_7 ,\custom_alu/mult/mult16_1/PSUM3__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_1/PSUM3__60_carry_n_4 ,\custom_alu/mult/mult16_1/PSUM3__60_carry_n_5 ,\custom_alu/mult/mult16_1/PSUM3__60_carry_n_6 ,\custom_alu/mult/mult16_1/PSUM3__60_carry_n_7 }),
        .S({PSUM3__60_carry_i_2__1_n_0,PSUM3__60_carry_i_3__1_n_0,PSUM3__60_carry_i_4__1_n_0,PSUM3__60_carry_i_5__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__60_carry__0 
       (.CI(\custom_alu/mult/mult16_1/PSUM3__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_0 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_1 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_2 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__0_i_1__1_n_0,PSUM3__60_carry__0_i_2__1_n_0,PSUM3__60_carry__0_i_3__1_n_0,PSUM3__60_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_4 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_5 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_6 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_7 }),
        .S({PSUM3__60_carry__0_i_5__1_n_0,PSUM3__60_carry__0_i_6__1_n_0,PSUM3__60_carry__0_i_7__1_n_0,PSUM3__60_carry__0_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__60_carry__1 
       (.CI(\custom_alu/mult/mult16_1/PSUM3__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_0 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_1 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_2 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__1_i_1__1_n_0,PSUM3__60_carry__1_i_2__2_n_0,PSUM3__60_carry__1_i_3__1_n_0,PSUM3__60_carry__1_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_4 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_5 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_6 ,\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_7 }),
        .S({PSUM3__60_carry__1_i_5__2_n_0,PSUM3__60_carry__1_i_6__2_n_0,PSUM3__60_carry__1_i_7__2_n_0,PSUM3__60_carry__1_i_8__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/PSUM3__60_carry__2 
       (.CI(\custom_alu/mult/mult16_1/PSUM3__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_1/PSUM3__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM3__60_carry__2_i_1__2_n_0}));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[11]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[43] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[27] ),
        .O(\custom_alu/mult/mult16_1/Q[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[11]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[42] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[26] ),
        .O(\custom_alu/mult/mult16_1/Q[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[11]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[25] ),
        .O(\custom_alu/mult/mult16_1/Q[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[11]_i_5 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[24] ),
        .O(\custom_alu/mult/mult16_1/Q[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[15]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[47] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[31] ),
        .O(\custom_alu/mult/mult16_1/Q[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[15]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[46] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[30] ),
        .O(\custom_alu/mult/mult16_1/Q[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[15]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[45] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[29] ),
        .O(\custom_alu/mult/mult16_1/Q[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[15]_i_5 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[44] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[28] ),
        .O(\custom_alu/mult/mult16_1/Q[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[3]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[19] ),
        .O(\custom_alu/mult/mult16_1/Q[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[3]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[18] ),
        .O(\custom_alu/mult/mult16_1/Q[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[3]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[17] ),
        .O(\custom_alu/mult/mult16_1/Q[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[3]_i_5 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/mult16_1/Q[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[74]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[27] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[2] ),
        .O(\custom_alu/mult/mult16_1/Q[74]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[74]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[26] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[1] ),
        .O(\custom_alu/mult/mult16_1/Q[74]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[74]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[25] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[0] ),
        .O(\custom_alu/mult/mult16_1/Q[74]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[78]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[31] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[6] ),
        .O(\custom_alu/mult/mult16_1/Q[78]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[78]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[30] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[5] ),
        .O(\custom_alu/mult/mult16_1/Q[78]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[78]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[29] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[4] ),
        .O(\custom_alu/mult/mult16_1/Q[78]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[78]_i_5 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[28] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[3] ),
        .O(\custom_alu/mult/mult16_1/Q[78]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[7]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[23] ),
        .O(\custom_alu/mult/mult16_1/Q[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[7]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[22] ),
        .O(\custom_alu/mult/mult16_1/Q[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[7]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[21] ),
        .O(\custom_alu/mult/mult16_1/Q[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[7]_i_5 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[20] ),
        .O(\custom_alu/mult/mult16_1/Q[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[82]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[10] ),
        .O(\custom_alu/mult/mult16_1/Q[82]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[82]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[9] ),
        .O(\custom_alu/mult/mult16_1/Q[82]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[82]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[8] ),
        .O(\custom_alu/mult/mult16_1/Q[82]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[82]_i_5 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[7] ),
        .O(\custom_alu/mult/mult16_1/Q[82]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[86]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[14] ),
        .O(\custom_alu/mult/mult16_1/Q[86]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[86]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[13] ),
        .O(\custom_alu/mult/mult16_1/Q[86]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[86]_i_4 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[12] ),
        .O(\custom_alu/mult/mult16_1/Q[86]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[86]_i_5 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[11] ),
        .O(\custom_alu/mult/mult16_1/Q[86]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[90]_i_2 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/mult16_1/Q[90]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_1/Q[90]_i_3 
       (.I0(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[15] ),
        .O(\custom_alu/mult/mult16_1/Q[90]_i_3_n_0 ));
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[11]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[43] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[42] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[41] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[40] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[11]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[11]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[11]_i_4_n_0 ,\custom_alu/mult/mult16_1/Q[11]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[15]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[11]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[47] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[46] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[45] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[44] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[15]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[15]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[15]_i_4_n_0 ,\custom_alu/mult/mult16_1/Q[15]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[16]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[15]_i_1_n_0 ),
        .CO(\custom_alu/mult/mult16_1/Q_reg[16]_i_1_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[35] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[34] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[33] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[32] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[3]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[3]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[3]_i_4_n_0 ,\custom_alu/mult/mult16_1/Q[3]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[74]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[27] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[26] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[25] ,\<const0> }),
        .O({\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[74]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[74]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[74]_i_4_n_0 ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[24] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[78]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[74]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[31] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[30] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[29] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[28] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[78]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[78]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[78]_i_4_n_0 ,\custom_alu/mult/mult16_1/Q[78]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[7]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[3]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[39] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[38] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[37] ,\custom_alu/mult/mult16_1/FF_MULT_0/Q_reg_n_0_[36] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[7]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[7]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[7]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[7]_i_4_n_0 ,\custom_alu/mult/mult16_1/Q[7]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[82]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[78]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[35] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[34] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[33] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[32] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[82]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[82]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[82]_i_4_n_0 ,\custom_alu/mult/mult16_1/Q[82]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[86]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[82]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[39] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[38] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[37] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[36] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/Q[86]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[86]_i_3_n_0 ,\custom_alu/mult/mult16_1/Q[86]_i_4_n_0 ,\custom_alu/mult/mult16_1/Q[86]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[90]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[86]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[41] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[40] }),
        .O({\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[43] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[42] ,\custom_alu/mult/mult16_1/Q[90]_i_2_n_0 ,\custom_alu/mult/mult16_1/Q[90]_i_3_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[94]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[90]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_0 ,\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_1 ,\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_2 ,\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_4 ,\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_5 ,\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_6 ,\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[47] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[46] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[45] ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[44] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_1/Q_reg[95]_i_1 
       (.CI(\custom_alu/mult/mult16_1/Q_reg[94]_i_1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_1/Q_reg[95]_i_1_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,\custom_alu/mult/mult16_1/FF_MULT_1/Q_reg_n_0_[48] }));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM2__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM1__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[49] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[49] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[50] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[50] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[51] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[51] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[52] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[52] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[53] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[53] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[54] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[54] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM0__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[63] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_0/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[9] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[16]_i_1_n_3 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[48] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[49] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[50] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[51] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[52] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[53] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[54] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[55] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[56] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[57] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[58] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[59] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[60] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[61] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[62] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[63] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[0] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[1] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[2] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[3] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[4] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[5] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[6] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[7] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[8] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[9] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[10] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[11] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[12] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[13] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[14] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[15] ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_2/FF_MULT_1/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[9] ),
        .R(RST0));
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__0_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM0__0_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM0__0_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM0__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry_i_1__0_n_0,PSUM0__0_carry_i_2__1_n_0,PSUM0__0_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM0__0_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM0__0_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM0__0_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM0__0_carry_n_7 }),
        .S({PSUM0__0_carry_i_4__1_n_0,PSUM0__0_carry_i_5__1_n_0,PSUM0__0_carry_i_6__0_n_0,PSUM0__0_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__0_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM0__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry__0_i_1__0_n_0,PSUM0__0_carry__0_i_2__0_n_0,PSUM0__0_carry__0_i_3__1_n_0,PSUM0__0_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_7 }),
        .S({PSUM0__0_carry__0_i_5__0_n_0,PSUM0__0_carry__0_i_6__0_n_0,PSUM0__0_carry__0_i_7__1_n_0,PSUM0__0_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__0_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM0__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__0_carry__1_i_1__0_n_0,PSUM0__0_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__0_carry__1_i_3__0_n_0,PSUM0__0_carry__1_i_4__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__30_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM0__30_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM0__30_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM0__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry_i_1__1_n_0,PSUM0__30_carry_i_2__0_n_0,PSUM0__30_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM0__30_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM0__30_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM0__30_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM0__30_carry_n_7 }),
        .S({PSUM0__30_carry_i_4__1_n_0,PSUM0__30_carry_i_5__0_n_0,PSUM0__30_carry_i_6__0_n_0,PSUM0__30_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__30_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM0__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry__0_i_1__0_n_0,PSUM0__30_carry__0_i_2__1_n_0,PSUM0__30_carry__0_i_3__0_n_0,PSUM0__30_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_7 }),
        .S({PSUM0__30_carry__0_i_5__1_n_0,PSUM0__30_carry__0_i_6__1_n_0,PSUM0__30_carry__0_i_7__1_n_0,PSUM0__30_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__30_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM0__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM0__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__30_carry__1_i_1__0_n_0,PSUM0__30_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM0__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__30_carry__1_i_3__0_n_0,PSUM0__30_carry__1_i_4__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__60_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM0__60_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM0__60_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM0__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry_i_1__0_n_0,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM0__0_carry__0_n_7 ,\custom_alu/mult/mult16_2/PSUM0__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_2/PSUM0__60_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM0__60_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM0__60_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM0__60_carry_n_7 }),
        .S({PSUM0__60_carry_i_2__0_n_0,PSUM0__60_carry_i_3__0_n_0,PSUM0__60_carry_i_4__0_n_0,PSUM0__60_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__60_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM0__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__0_i_1__0_n_0,PSUM0__60_carry__0_i_2__0_n_0,PSUM0__60_carry__0_i_3__0_n_0,PSUM0__60_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_7 }),
        .S({PSUM0__60_carry__0_i_5__0_n_0,PSUM0__60_carry__0_i_6__0_n_0,PSUM0__60_carry__0_i_7__0_n_0,PSUM0__60_carry__0_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__60_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM0__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_0 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_1 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_2 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__1_i_1__0_n_0,PSUM0__60_carry__1_i_2__1_n_0,PSUM0__60_carry__1_i_3__0_n_0,PSUM0__60_carry__1_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_4 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_5 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_7 }),
        .S({PSUM0__60_carry__1_i_5__1_n_0,PSUM0__60_carry__1_i_6__1_n_0,PSUM0__60_carry__1_i_7__1_n_0,PSUM0__60_carry__1_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM0__60_carry__2 
       (.CI(\custom_alu/mult/mult16_2/PSUM0__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_2/PSUM0__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM0__60_carry__2_i_1__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__0_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM1__0_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM1__0_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM1__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry_i_1__0_n_0,PSUM1__0_carry_i_2__0_n_0,PSUM1__0_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM1__0_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM1__0_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM1__0_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM1__0_carry_n_7 }),
        .S({PSUM1__0_carry_i_4__0_n_0,PSUM1__0_carry_i_5__0_n_0,PSUM1__0_carry_i_6__0_n_0,PSUM1__0_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__0_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM1__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry__0_i_1__0_n_0,PSUM1__0_carry__0_i_2__0_n_0,PSUM1__0_carry__0_i_3__0_n_0,PSUM1__0_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_7 }),
        .S({PSUM1__0_carry__0_i_5__0_n_0,PSUM1__0_carry__0_i_6__0_n_0,PSUM1__0_carry__0_i_7__0_n_0,PSUM1__0_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__0_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM1__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__0_carry__1_i_1__0_n_0,PSUM1__0_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__0_carry__1_i_3__0_n_0,PSUM1__0_carry__1_i_4__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__30_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM1__30_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM1__30_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM1__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry_i_1__0_n_0,PSUM1__30_carry_i_2__0_n_0,PSUM1__30_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM1__30_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM1__30_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM1__30_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM1__30_carry_n_7 }),
        .S({PSUM1__30_carry_i_4__0_n_0,PSUM1__30_carry_i_5__0_n_0,PSUM1__30_carry_i_6__0_n_0,PSUM1__30_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__30_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM1__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry__0_i_1__0_n_0,PSUM1__30_carry__0_i_2__0_n_0,PSUM1__30_carry__0_i_3__0_n_0,PSUM1__30_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_7 }),
        .S({PSUM1__30_carry__0_i_5__0_n_0,PSUM1__30_carry__0_i_6__0_n_0,PSUM1__30_carry__0_i_7__0_n_0,PSUM1__30_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__30_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM1__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM1__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__30_carry__1_i_1__0_n_0,PSUM1__30_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM1__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__30_carry__1_i_3__0_n_0,PSUM1__30_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__60_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM1__60_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM1__60_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM1__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry_i_1__0_n_0,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM1__0_carry__0_n_7 ,\custom_alu/mult/mult16_2/PSUM1__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_2/PSUM1__60_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM1__60_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM1__60_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM1__60_carry_n_7 }),
        .S({PSUM1__60_carry_i_2__0_n_0,PSUM1__60_carry_i_3__0_n_0,PSUM1__60_carry_i_4__0_n_0,PSUM1__60_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__60_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM1__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__0_i_1__0_n_0,PSUM1__60_carry__0_i_2__0_n_0,PSUM1__60_carry__0_i_3__0_n_0,PSUM1__60_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_7 }),
        .S({PSUM1__60_carry__0_i_5__0_n_0,PSUM1__60_carry__0_i_6__0_n_0,PSUM1__60_carry__0_i_7__0_n_0,PSUM1__60_carry__0_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__60_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM1__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_0 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_1 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_2 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__1_i_1__0_n_0,PSUM1__60_carry__1_i_2__0_n_0,PSUM1__60_carry__1_i_3__0_n_0,PSUM1__60_carry__1_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_4 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_5 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_7 }),
        .S({PSUM1__60_carry__1_i_5__0_n_0,PSUM1__60_carry__1_i_6__0_n_0,PSUM1__60_carry__1_i_7__0_n_0,PSUM1__60_carry__1_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM1__60_carry__2 
       (.CI(\custom_alu/mult/mult16_2/PSUM1__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_2/PSUM1__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM1__60_carry__2_i_1__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__0_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM2__0_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM2__0_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM2__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry_i_1__0_n_0,PSUM2__0_carry_i_2__0_n_0,PSUM2__0_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM2__0_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM2__0_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM2__0_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM2__0_carry_n_7 }),
        .S({PSUM2__0_carry_i_4__0_n_0,PSUM2__0_carry_i_5__0_n_0,PSUM2__0_carry_i_6__0_n_0,PSUM2__0_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__0_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM2__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry__0_i_1__0_n_0,PSUM2__0_carry__0_i_2__0_n_0,PSUM2__0_carry__0_i_3__0_n_0,PSUM2__0_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_7 }),
        .S({PSUM2__0_carry__0_i_5__0_n_0,PSUM2__0_carry__0_i_6__0_n_0,PSUM2__0_carry__0_i_7__0_n_0,PSUM2__0_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__0_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM2__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__0_carry__1_i_1__0_n_0,PSUM2__0_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__0_carry__1_i_3__0_n_0,PSUM2__0_carry__1_i_4__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__30_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM2__30_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM2__30_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM2__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry_i_1__0_n_0,PSUM2__30_carry_i_2__0_n_0,PSUM2__30_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM2__30_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM2__30_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM2__30_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM2__30_carry_n_7 }),
        .S({PSUM2__30_carry_i_4__0_n_0,PSUM2__30_carry_i_5__0_n_0,PSUM2__30_carry_i_6__0_n_0,PSUM2__30_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__30_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM2__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry__0_i_1__0_n_0,PSUM2__30_carry__0_i_2__0_n_0,PSUM2__30_carry__0_i_3__0_n_0,PSUM2__30_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_7 }),
        .S({PSUM2__30_carry__0_i_5__0_n_0,PSUM2__30_carry__0_i_6__0_n_0,PSUM2__30_carry__0_i_7__0_n_0,PSUM2__30_carry__0_i_8__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__30_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM2__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM2__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__30_carry__1_i_1__0_n_0,PSUM2__30_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM2__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__30_carry__1_i_3__0_n_0,PSUM2__30_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__60_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM2__60_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM2__60_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM2__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry_i_1__0_n_0,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM2__0_carry__0_n_7 ,\custom_alu/mult/mult16_2/PSUM2__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_2/PSUM2__60_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM2__60_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM2__60_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM2__60_carry_n_7 }),
        .S({PSUM2__60_carry_i_2__0_n_0,PSUM2__60_carry_i_3__0_n_0,PSUM2__60_carry_i_4__0_n_0,PSUM2__60_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__60_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM2__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__0_i_1__0_n_0,PSUM2__60_carry__0_i_2__0_n_0,PSUM2__60_carry__0_i_3__0_n_0,PSUM2__60_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_7 }),
        .S({PSUM2__60_carry__0_i_5__0_n_0,PSUM2__60_carry__0_i_6__0_n_0,PSUM2__60_carry__0_i_7__0_n_0,PSUM2__60_carry__0_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__60_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM2__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_0 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_1 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_2 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__1_i_1__0_n_0,PSUM2__60_carry__1_i_2__0_n_0,PSUM2__60_carry__1_i_3__0_n_0,PSUM2__60_carry__1_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_4 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_5 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_7 }),
        .S({PSUM2__60_carry__1_i_5__0_n_0,PSUM2__60_carry__1_i_6__0_n_0,PSUM2__60_carry__1_i_7__0_n_0,PSUM2__60_carry__1_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM2__60_carry__2 
       (.CI(\custom_alu/mult/mult16_2/PSUM2__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_2/PSUM2__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM2__60_carry__2_i_1__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__0_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM3__0_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM3__0_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM3__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry_i_1__0_n_0,PSUM3__0_carry_i_2__1_n_0,PSUM3__0_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM3__0_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM3__0_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM3__0_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM3__0_carry_n_7 }),
        .S({PSUM3__0_carry_i_4__1_n_0,PSUM3__0_carry_i_5__1_n_0,PSUM3__0_carry_i_6__0_n_0,PSUM3__0_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__0_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM3__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry__0_i_1__0_n_0,PSUM3__0_carry__0_i_2__0_n_0,PSUM3__0_carry__0_i_3__1_n_0,PSUM3__0_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_7 }),
        .S({PSUM3__0_carry__0_i_5__0_n_0,PSUM3__0_carry__0_i_6__0_n_0,PSUM3__0_carry__0_i_7__1_n_0,PSUM3__0_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__0_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM3__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__0_carry__1_i_1__0_n_0,PSUM3__0_carry__1_i_2__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__0_carry__1_i_3__0_n_0,PSUM3__0_carry__1_i_4__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__30_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM3__30_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM3__30_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM3__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry_i_1__1_n_0,PSUM3__30_carry_i_2__0_n_0,PSUM3__30_carry_i_3__0_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_2/PSUM3__30_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM3__30_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM3__30_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM3__30_carry_n_7 }),
        .S({PSUM3__30_carry_i_4__1_n_0,PSUM3__30_carry_i_5__0_n_0,PSUM3__30_carry_i_6__0_n_0,PSUM3__30_carry_i_7__2_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__30_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM3__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry__0_i_1__0_n_0,PSUM3__30_carry__0_i_2__1_n_0,PSUM3__30_carry__0_i_3__0_n_0,PSUM3__30_carry__0_i_4__1_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_7 }),
        .S({PSUM3__30_carry__0_i_5__1_n_0,PSUM3__30_carry__0_i_6__1_n_0,PSUM3__30_carry__0_i_7__1_n_0,PSUM3__30_carry__0_i_8__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__30_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM3__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_2/PSUM3__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__30_carry__1_i_1__0_n_0,PSUM3__30_carry__1_i_2__1_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM3__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__30_carry__1_i_3__0_n_0,PSUM3__30_carry__1_i_4__1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__60_carry_n_0 ,\custom_alu/mult/mult16_2/PSUM3__60_carry_n_1 ,\custom_alu/mult/mult16_2/PSUM3__60_carry_n_2 ,\custom_alu/mult/mult16_2/PSUM3__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry_i_1__0_n_0,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM3__0_carry__0_n_7 ,\custom_alu/mult/mult16_2/PSUM3__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_2/PSUM3__60_carry_n_4 ,\custom_alu/mult/mult16_2/PSUM3__60_carry_n_5 ,\custom_alu/mult/mult16_2/PSUM3__60_carry_n_6 ,\custom_alu/mult/mult16_2/PSUM3__60_carry_n_7 }),
        .S({PSUM3__60_carry_i_2__0_n_0,PSUM3__60_carry_i_3__0_n_0,PSUM3__60_carry_i_4__0_n_0,PSUM3__60_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__60_carry__0 
       (.CI(\custom_alu/mult/mult16_2/PSUM3__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_0 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_1 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_2 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__0_i_1__0_n_0,PSUM3__60_carry__0_i_2__0_n_0,PSUM3__60_carry__0_i_3__0_n_0,PSUM3__60_carry__0_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_4 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_5 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_6 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_7 }),
        .S({PSUM3__60_carry__0_i_5__0_n_0,PSUM3__60_carry__0_i_6__0_n_0,PSUM3__60_carry__0_i_7__0_n_0,PSUM3__60_carry__0_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__60_carry__1 
       (.CI(\custom_alu/mult/mult16_2/PSUM3__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_0 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_1 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_2 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__1_i_1__0_n_0,PSUM3__60_carry__1_i_2__1_n_0,PSUM3__60_carry__1_i_3__0_n_0,PSUM3__60_carry__1_i_4__0_n_0}),
        .O({\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_4 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_5 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_6 ,\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_7 }),
        .S({PSUM3__60_carry__1_i_5__1_n_0,PSUM3__60_carry__1_i_6__1_n_0,PSUM3__60_carry__1_i_7__1_n_0,PSUM3__60_carry__1_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/PSUM3__60_carry__2 
       (.CI(\custom_alu/mult/mult16_2/PSUM3__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_2/PSUM3__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM3__60_carry__2_i_1__1_n_0}));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[11]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[43] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[27] ),
        .O(\custom_alu/mult/mult16_2/Q[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[11]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[42] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[26] ),
        .O(\custom_alu/mult/mult16_2/Q[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[11]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[25] ),
        .O(\custom_alu/mult/mult16_2/Q[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[11]_i_5 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[24] ),
        .O(\custom_alu/mult/mult16_2/Q[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[15]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[47] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[31] ),
        .O(\custom_alu/mult/mult16_2/Q[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[15]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[46] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[30] ),
        .O(\custom_alu/mult/mult16_2/Q[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[15]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[45] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[29] ),
        .O(\custom_alu/mult/mult16_2/Q[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[15]_i_5 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[44] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[28] ),
        .O(\custom_alu/mult/mult16_2/Q[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[3]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[19] ),
        .O(\custom_alu/mult/mult16_2/Q[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[3]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[18] ),
        .O(\custom_alu/mult/mult16_2/Q[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[3]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[17] ),
        .O(\custom_alu/mult/mult16_2/Q[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[3]_i_5 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/mult16_2/Q[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[42]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[27] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[2] ),
        .O(\custom_alu/mult/mult16_2/Q[42]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[42]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[26] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[1] ),
        .O(\custom_alu/mult/mult16_2/Q[42]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[42]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[25] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[0] ),
        .O(\custom_alu/mult/mult16_2/Q[42]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[46]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[31] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[6] ),
        .O(\custom_alu/mult/mult16_2/Q[46]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[46]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[30] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[5] ),
        .O(\custom_alu/mult/mult16_2/Q[46]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[46]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[29] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[4] ),
        .O(\custom_alu/mult/mult16_2/Q[46]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[46]_i_5 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[28] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[3] ),
        .O(\custom_alu/mult/mult16_2/Q[46]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[50]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[10] ),
        .O(\custom_alu/mult/mult16_2/Q[50]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[50]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[9] ),
        .O(\custom_alu/mult/mult16_2/Q[50]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[50]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[8] ),
        .O(\custom_alu/mult/mult16_2/Q[50]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[50]_i_5 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[7] ),
        .O(\custom_alu/mult/mult16_2/Q[50]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[54]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[14] ),
        .O(\custom_alu/mult/mult16_2/Q[54]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[54]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[13] ),
        .O(\custom_alu/mult/mult16_2/Q[54]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[54]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[12] ),
        .O(\custom_alu/mult/mult16_2/Q[54]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[54]_i_5 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[11] ),
        .O(\custom_alu/mult/mult16_2/Q[54]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[58]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/mult16_2/Q[58]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[58]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[15] ),
        .O(\custom_alu/mult/mult16_2/Q[58]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[7]_i_2 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[23] ),
        .O(\custom_alu/mult/mult16_2/Q[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[7]_i_3 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[22] ),
        .O(\custom_alu/mult/mult16_2/Q[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[7]_i_4 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[21] ),
        .O(\custom_alu/mult/mult16_2/Q[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_2/Q[7]_i_5 
       (.I0(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[20] ),
        .O(\custom_alu/mult/mult16_2/Q[7]_i_5_n_0 ));
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[11]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[43] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[42] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[41] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[40] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[11]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[11]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[11]_i_4_n_0 ,\custom_alu/mult/mult16_2/Q[11]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[15]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[11]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[47] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[46] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[45] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[44] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[15]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[15]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[15]_i_4_n_0 ,\custom_alu/mult/mult16_2/Q[15]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[16]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[15]_i_1_n_0 ),
        .CO(\custom_alu/mult/mult16_2/Q_reg[16]_i_1_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[35] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[34] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[33] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[32] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[3]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[3]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[3]_i_4_n_0 ,\custom_alu/mult/mult16_2/Q[3]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[42]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[27] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[26] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[25] ,\<const0> }),
        .O({\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[42]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[42]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[42]_i_4_n_0 ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[24] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[46]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[42]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[31] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[30] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[29] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[28] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[46]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[46]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[46]_i_4_n_0 ,\custom_alu/mult/mult16_2/Q[46]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[50]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[46]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[35] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[34] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[33] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[32] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[50]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[50]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[50]_i_4_n_0 ,\custom_alu/mult/mult16_2/Q[50]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[54]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[50]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[39] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[38] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[37] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[36] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[54]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[54]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[54]_i_4_n_0 ,\custom_alu/mult/mult16_2/Q[54]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[58]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[54]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[41] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[40] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[43] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[42] ,\custom_alu/mult/mult16_2/Q[58]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[58]_i_3_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[62]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[58]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[47] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[46] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[45] ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[44] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[63]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[62]_i_1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_2/Q_reg[63]_i_1_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,\custom_alu/mult/mult16_2/FF_MULT_1/Q_reg_n_0_[48] }));
  CARRY4 \custom_alu/mult/mult16_2/Q_reg[7]_i_1 
       (.CI(\custom_alu/mult/mult16_2/Q_reg[3]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_0 ,\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_1 ,\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_2 ,\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[39] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[38] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[37] ,\custom_alu/mult/mult16_2/FF_MULT_0/Q_reg_n_0_[36] }),
        .O({\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_4 ,\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_5 ,\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_6 ,\custom_alu/mult/mult16_2/Q_reg[7]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_2/Q[7]_i_2_n_0 ,\custom_alu/mult/mult16_2/Q[7]_i_3_n_0 ,\custom_alu/mult/mult16_2/Q[7]_i_4_n_0 ,\custom_alu/mult/mult16_2/Q[7]_i_5_n_0 }));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[16] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[17] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[17] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[18] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[18] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[19] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[19] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[1] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[20] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[20] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[21] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[21] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[22] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[22] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[23] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[23] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM2__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM1__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[55] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[55] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[56] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[56] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[57] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[57] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[58] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[58] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[59] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[59] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[60] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[60] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[61] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[61] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[62] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[62] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[63] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry__2_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[63] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[9] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\<const1> ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_r_n_0 ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[0] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[0] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[10] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[10] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[11] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[11] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[12] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[12] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[13] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[13] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[14] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[14] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[15] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[15] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[16] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[16]_i_1_n_3 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[16] ),
        .R(RST0));
  (* srl_bus_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/mult16_3/PSUM0__0_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[17]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/mult16_3/PSUM0__0_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[18]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/mult16_3/PSUM0__0_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[19]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[1] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[1] ),
        .R(RST0));
  (* srl_bus_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[20]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[21]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[22]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  (* srl_bus_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg " *) 
  (* srl_name = "\\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r 
       (.A0(\<const1> ),
        .A1(\<const0> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(CLK_IBUF_BUFG),
        .D(\custom_alu/mult/mult16_3/PSUM0__60_carry_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[23]_srl2___custom_alu_mult_mult16_3_FF_MULT_1_Q_reg_r_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[24] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[55] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[24] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[25] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[56] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[25] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[26] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[57] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[26] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[27] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[58] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[27] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[28] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[59] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[28] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[29] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[60] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[29] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[2] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[2] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[30] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[61] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[30] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[31] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[62] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[31] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[32] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[63] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[32] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[33] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[0] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[33] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[34] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[1] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[34] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[35] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[2] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[35] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[36] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[3] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[36] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[37] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[4] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[37] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[38] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[5] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[38] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[39] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[6] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[39] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[3] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[3] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[40] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[7] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[40] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[41] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[8] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[41] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[42] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[9] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[42] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[43] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[10] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[43] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[44] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[11] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[44] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[45] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[12] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[45] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[46] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[13] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[46] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[47] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[14] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[47] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[48] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[15] ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[48] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[4] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[4] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[5] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[5] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[6] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_5 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[6] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[7] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_4 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[7] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[8] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_7 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[8] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg[9] 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_6 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[9] ),
        .R(RST0));
  FDRE #(
    .INIT(1'b0)) 
    \custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_r 
       (.C(CLK_IBUF_BUFG),
        .CE(\<const1> ),
        .D(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_r_n_0 ),
        .Q(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_r_n_0 ),
        .R(RST0));
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__0_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM0__0_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM0__0_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM0__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry_i_1_n_0,PSUM0__0_carry_i_2_n_0,PSUM0__0_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM0__0_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM0__0_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM0__0_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM0__0_carry_n_7 }),
        .S({PSUM0__0_carry_i_4_n_0,PSUM0__0_carry_i_5_n_0,PSUM0__0_carry_i_6_n_0,PSUM0__0_carry_i_7__1_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__0_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM0__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__0_carry__0_i_1_n_0,PSUM0__0_carry__0_i_2_n_0,PSUM0__0_carry__0_i_3_n_0,PSUM0__0_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_7 }),
        .S({PSUM0__0_carry__0_i_5_n_0,PSUM0__0_carry__0_i_6_n_0,PSUM0__0_carry__0_i_7_n_0,PSUM0__0_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__0_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM0__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__0_carry__1_i_1_n_0,PSUM0__0_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__0_carry__1_i_3_n_0,PSUM0__0_carry__1_i_4_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__30_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM0__30_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM0__30_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM0__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry_i_1_n_0,PSUM0__30_carry_i_2_n_0,PSUM0__30_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM0__30_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM0__30_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM0__30_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM0__30_carry_n_7 }),
        .S({PSUM0__30_carry_i_4_n_0,PSUM0__30_carry_i_5_n_0,PSUM0__30_carry_i_6_n_0,PSUM0__30_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__30_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM0__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__30_carry__0_i_1_n_0,PSUM0__30_carry__0_i_2__0_n_0,PSUM0__30_carry__0_i_3_n_0,PSUM0__30_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_7 }),
        .S({PSUM0__30_carry__0_i_5_n_0,PSUM0__30_carry__0_i_6__0_n_0,PSUM0__30_carry__0_i_7__0_n_0,PSUM0__30_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__30_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM0__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM0__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM0__30_carry__1_i_1_n_0,PSUM0__30_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM0__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM0__30_carry__1_i_3_n_0,PSUM0__30_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__60_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM0__60_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM0__60_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM0__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry_i_1_n_0,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM0__0_carry__0_n_7 ,\custom_alu/mult/mult16_3/PSUM0__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_3/PSUM0__60_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM0__60_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM0__60_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM0__60_carry_n_7 }),
        .S({PSUM0__60_carry_i_2_n_0,PSUM0__60_carry_i_3_n_0,PSUM0__60_carry_i_4_n_0,PSUM0__60_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__60_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM0__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__0_i_1_n_0,PSUM0__60_carry__0_i_2_n_0,PSUM0__60_carry__0_i_3_n_0,PSUM0__60_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_7 }),
        .S({PSUM0__60_carry__0_i_5_n_0,PSUM0__60_carry__0_i_6_n_0,PSUM0__60_carry__0_i_7_n_0,PSUM0__60_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__60_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM0__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_0 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_1 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_2 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM0__60_carry__1_i_1_n_0,PSUM0__60_carry__1_i_2_n_0,PSUM0__60_carry__1_i_3_n_0,PSUM0__60_carry__1_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_4 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_5 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_7 }),
        .S({PSUM0__60_carry__1_i_5_n_0,PSUM0__60_carry__1_i_6_n_0,PSUM0__60_carry__1_i_7_n_0,PSUM0__60_carry__1_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM0__60_carry__2 
       (.CI(\custom_alu/mult/mult16_3/PSUM0__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_3/PSUM0__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM0__60_carry__2_i_1_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__0_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM1__0_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM1__0_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM1__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry_i_1_n_0,PSUM1__0_carry_i_2_n_0,PSUM1__0_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM1__0_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM1__0_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM1__0_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM1__0_carry_n_7 }),
        .S({PSUM1__0_carry_i_4_n_0,PSUM1__0_carry_i_5_n_0,PSUM1__0_carry_i_6_n_0,PSUM1__0_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__0_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM1__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__0_carry__0_i_1_n_0,PSUM1__0_carry__0_i_2_n_0,PSUM1__0_carry__0_i_3_n_0,PSUM1__0_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_7 }),
        .S({PSUM1__0_carry__0_i_5_n_0,PSUM1__0_carry__0_i_6_n_0,PSUM1__0_carry__0_i_7_n_0,PSUM1__0_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__0_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM1__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__0_carry__1_i_1_n_0,PSUM1__0_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__0_carry__1_i_3_n_0,PSUM1__0_carry__1_i_4_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__30_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM1__30_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM1__30_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM1__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry_i_1_n_0,PSUM1__30_carry_i_2_n_0,PSUM1__30_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM1__30_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM1__30_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM1__30_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM1__30_carry_n_7 }),
        .S({PSUM1__30_carry_i_4_n_0,PSUM1__30_carry_i_5_n_0,PSUM1__30_carry_i_6_n_0,PSUM1__30_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__30_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM1__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__30_carry__0_i_1_n_0,PSUM1__30_carry__0_i_2_n_0,PSUM1__30_carry__0_i_3_n_0,PSUM1__30_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_7 }),
        .S({PSUM1__30_carry__0_i_5_n_0,PSUM1__30_carry__0_i_6_n_0,PSUM1__30_carry__0_i_7_n_0,PSUM1__30_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__30_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM1__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM1__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM1__30_carry__1_i_1_n_0,PSUM1__30_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM1__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM1__30_carry__1_i_3_n_0,PSUM1__30_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__60_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM1__60_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM1__60_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM1__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry_i_1_n_0,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM1__0_carry__0_n_7 ,\custom_alu/mult/mult16_3/PSUM1__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_3/PSUM1__60_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM1__60_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM1__60_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM1__60_carry_n_7 }),
        .S({PSUM1__60_carry_i_2_n_0,PSUM1__60_carry_i_3_n_0,PSUM1__60_carry_i_4_n_0,PSUM1__60_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__60_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM1__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__0_i_1_n_0,PSUM1__60_carry__0_i_2_n_0,PSUM1__60_carry__0_i_3_n_0,PSUM1__60_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_7 }),
        .S({PSUM1__60_carry__0_i_5_n_0,PSUM1__60_carry__0_i_6_n_0,PSUM1__60_carry__0_i_7_n_0,PSUM1__60_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__60_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM1__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_0 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_1 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_2 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM1__60_carry__1_i_1_n_0,PSUM1__60_carry__1_i_2_n_0,PSUM1__60_carry__1_i_3_n_0,PSUM1__60_carry__1_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_4 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_5 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_7 }),
        .S({PSUM1__60_carry__1_i_5_n_0,PSUM1__60_carry__1_i_6_n_0,PSUM1__60_carry__1_i_7_n_0,PSUM1__60_carry__1_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM1__60_carry__2 
       (.CI(\custom_alu/mult/mult16_3/PSUM1__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_3/PSUM1__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM1__60_carry__2_i_1_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__0_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM2__0_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM2__0_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM2__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry_i_1_n_0,PSUM2__0_carry_i_2_n_0,PSUM2__0_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM2__0_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM2__0_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM2__0_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM2__0_carry_n_7 }),
        .S({PSUM2__0_carry_i_4_n_0,PSUM2__0_carry_i_5_n_0,PSUM2__0_carry_i_6_n_0,PSUM2__0_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__0_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM2__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__0_carry__0_i_1_n_0,PSUM2__0_carry__0_i_2_n_0,PSUM2__0_carry__0_i_3_n_0,PSUM2__0_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_7 }),
        .S({PSUM2__0_carry__0_i_5_n_0,PSUM2__0_carry__0_i_6_n_0,PSUM2__0_carry__0_i_7_n_0,PSUM2__0_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__0_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM2__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__0_carry__1_i_1_n_0,PSUM2__0_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__0_carry__1_i_3_n_0,PSUM2__0_carry__1_i_4_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__30_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM2__30_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM2__30_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM2__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry_i_1_n_0,PSUM2__30_carry_i_2_n_0,PSUM2__30_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM2__30_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM2__30_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM2__30_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM2__30_carry_n_7 }),
        .S({PSUM2__30_carry_i_4_n_0,PSUM2__30_carry_i_5_n_0,PSUM2__30_carry_i_6_n_0,PSUM2__30_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__30_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM2__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__30_carry__0_i_1_n_0,PSUM2__30_carry__0_i_2_n_0,PSUM2__30_carry__0_i_3_n_0,PSUM2__30_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_7 }),
        .S({PSUM2__30_carry__0_i_5_n_0,PSUM2__30_carry__0_i_6_n_0,PSUM2__30_carry__0_i_7_n_0,PSUM2__30_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__30_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM2__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM2__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM2__30_carry__1_i_1_n_0,PSUM2__30_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM2__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM2__30_carry__1_i_3_n_0,PSUM2__30_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__60_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM2__60_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM2__60_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM2__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry_i_1_n_0,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM2__0_carry__0_n_7 ,\custom_alu/mult/mult16_3/PSUM2__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_3/PSUM2__60_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM2__60_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM2__60_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM2__60_carry_n_7 }),
        .S({PSUM2__60_carry_i_2_n_0,PSUM2__60_carry_i_3_n_0,PSUM2__60_carry_i_4_n_0,PSUM2__60_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__60_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM2__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__0_i_1_n_0,PSUM2__60_carry__0_i_2_n_0,PSUM2__60_carry__0_i_3_n_0,PSUM2__60_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_7 }),
        .S({PSUM2__60_carry__0_i_5_n_0,PSUM2__60_carry__0_i_6_n_0,PSUM2__60_carry__0_i_7_n_0,PSUM2__60_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__60_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM2__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_0 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_1 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_2 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM2__60_carry__1_i_1_n_0,PSUM2__60_carry__1_i_2_n_0,PSUM2__60_carry__1_i_3_n_0,PSUM2__60_carry__1_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_4 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_5 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_7 }),
        .S({PSUM2__60_carry__1_i_5_n_0,PSUM2__60_carry__1_i_6_n_0,PSUM2__60_carry__1_i_7_n_0,PSUM2__60_carry__1_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM2__60_carry__2 
       (.CI(\custom_alu/mult/mult16_3/PSUM2__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_3/PSUM2__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM2__60_carry__2_i_1_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__0_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__0_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM3__0_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM3__0_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM3__0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry_i_1_n_0,PSUM3__0_carry_i_2_n_0,PSUM3__0_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM3__0_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM3__0_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM3__0_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM3__0_carry_n_7 }),
        .S({PSUM3__0_carry_i_4_n_0,PSUM3__0_carry_i_5_n_0,PSUM3__0_carry_i_6_n_0,PSUM3__0_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__0_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM3__0_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__0_carry__0_i_1_n_0,PSUM3__0_carry__0_i_2_n_0,PSUM3__0_carry__0_i_3_n_0,PSUM3__0_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_7 }),
        .S({PSUM3__0_carry__0_i_5_n_0,PSUM3__0_carry__0_i_6_n_0,PSUM3__0_carry__0_i_7_n_0,PSUM3__0_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__0_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM3__0_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__0_carry__1_i_1_n_0,PSUM3__0_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__0_carry__1_i_3_n_0,PSUM3__0_carry__1_i_4_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__30_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__30_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM3__30_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM3__30_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM3__30_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry_i_1_n_0,PSUM3__30_carry_i_2_n_0,PSUM3__30_carry_i_3_n_0,\<const0> }),
        .O({\custom_alu/mult/mult16_3/PSUM3__30_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM3__30_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM3__30_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM3__30_carry_n_7 }),
        .S({PSUM3__30_carry_i_4_n_0,PSUM3__30_carry_i_5_n_0,PSUM3__30_carry_i_6_n_0,PSUM3__30_carry_i_7__0_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__30_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM3__30_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__30_carry__0_i_1_n_0,PSUM3__30_carry__0_i_2_n_0,PSUM3__30_carry__0_i_3_n_0,PSUM3__30_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_7 }),
        .S({PSUM3__30_carry__0_i_5_n_0,PSUM3__30_carry__0_i_6_n_0,PSUM3__30_carry__0_i_7_n_0,PSUM3__30_carry__0_i_8_n_0}));
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__30_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM3__30_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_1 ,\NLW_custom_alu/mult/mult16_3/PSUM3__30_carry__1_CO_UNCONNECTED [1],\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,PSUM3__30_carry__1_i_1_n_0,PSUM3__30_carry__1_i_2_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM3__30_carry__1_n_7 }),
        .S({\<const0> ,\<const1> ,PSUM3__30_carry__1_i_3_n_0,PSUM3__30_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__60_carry 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__60_carry_n_0 ,\custom_alu/mult/mult16_3/PSUM3__60_carry_n_1 ,\custom_alu/mult/mult16_3/PSUM3__60_carry_n_2 ,\custom_alu/mult/mult16_3/PSUM3__60_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry_i_1_n_0,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM3__0_carry__0_n_7 ,\custom_alu/mult/mult16_3/PSUM3__0_carry_n_4 }),
        .O({\custom_alu/mult/mult16_3/PSUM3__60_carry_n_4 ,\custom_alu/mult/mult16_3/PSUM3__60_carry_n_5 ,\custom_alu/mult/mult16_3/PSUM3__60_carry_n_6 ,\custom_alu/mult/mult16_3/PSUM3__60_carry_n_7 }),
        .S({PSUM3__60_carry_i_2_n_0,PSUM3__60_carry_i_3_n_0,PSUM3__60_carry_i_4_n_0,PSUM3__60_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__60_carry__0 
       (.CI(\custom_alu/mult/mult16_3/PSUM3__60_carry_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_0 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_1 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_2 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__0_i_1_n_0,PSUM3__60_carry__0_i_2_n_0,PSUM3__60_carry__0_i_3_n_0,PSUM3__60_carry__0_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_4 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_5 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_6 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_7 }),
        .S({PSUM3__60_carry__0_i_5_n_0,PSUM3__60_carry__0_i_6_n_0,PSUM3__60_carry__0_i_7_n_0,PSUM3__60_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__60_carry__1 
       (.CI(\custom_alu/mult/mult16_3/PSUM3__60_carry__0_n_0 ),
        .CO({\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_0 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_1 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_2 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({PSUM3__60_carry__1_i_1_n_0,PSUM3__60_carry__1_i_2_n_0,PSUM3__60_carry__1_i_3_n_0,PSUM3__60_carry__1_i_4_n_0}),
        .O({\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_4 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_5 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_6 ,\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_7 }),
        .S({PSUM3__60_carry__1_i_5_n_0,PSUM3__60_carry__1_i_6_n_0,PSUM3__60_carry__1_i_7_n_0,PSUM3__60_carry__1_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/PSUM3__60_carry__2 
       (.CI(\custom_alu/mult/mult16_3/PSUM3__60_carry__1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_3/PSUM3__60_carry__2_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,PSUM3__60_carry__2_i_1_n_0}));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[10]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[27] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[2] ),
        .O(\custom_alu/mult/mult16_3/Q[10]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[10]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[26] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[1] ),
        .O(\custom_alu/mult/mult16_3/Q[10]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[10]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[25] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[0] ),
        .O(\custom_alu/mult/mult16_3/Q[10]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[11]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[43] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[27] ),
        .O(\custom_alu/mult/mult16_3/Q[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[11]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[42] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[26] ),
        .O(\custom_alu/mult/mult16_3/Q[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[11]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[25] ),
        .O(\custom_alu/mult/mult16_3/Q[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[11]_i_5 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[24] ),
        .O(\custom_alu/mult/mult16_3/Q[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[14]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[31] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[6] ),
        .O(\custom_alu/mult/mult16_3/Q[14]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[14]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[30] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[5] ),
        .O(\custom_alu/mult/mult16_3/Q[14]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[14]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[29] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[4] ),
        .O(\custom_alu/mult/mult16_3/Q[14]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[14]_i_5 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[28] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[3] ),
        .O(\custom_alu/mult/mult16_3/Q[14]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[15]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[47] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[31] ),
        .O(\custom_alu/mult/mult16_3/Q[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[15]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[46] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[30] ),
        .O(\custom_alu/mult/mult16_3/Q[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[15]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[45] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[29] ),
        .O(\custom_alu/mult/mult16_3/Q[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[15]_i_5 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[44] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[28] ),
        .O(\custom_alu/mult/mult16_3/Q[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[18]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[10] ),
        .O(\custom_alu/mult/mult16_3/Q[18]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[18]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[9] ),
        .O(\custom_alu/mult/mult16_3/Q[18]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[18]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[8] ),
        .O(\custom_alu/mult/mult16_3/Q[18]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[18]_i_5 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[7] ),
        .O(\custom_alu/mult/mult16_3/Q[18]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[22]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[14] ),
        .O(\custom_alu/mult/mult16_3/Q[22]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[22]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[13] ),
        .O(\custom_alu/mult/mult16_3/Q[22]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[22]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[12] ),
        .O(\custom_alu/mult/mult16_3/Q[22]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[22]_i_5 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[11] ),
        .O(\custom_alu/mult/mult16_3/Q[22]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[26]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[41] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/mult16_3/Q[26]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[26]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[40] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[15] ),
        .O(\custom_alu/mult/mult16_3/Q[26]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[3]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[35] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[19] ),
        .O(\custom_alu/mult/mult16_3/Q[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[3]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[34] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[18] ),
        .O(\custom_alu/mult/mult16_3/Q[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[3]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[33] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[17] ),
        .O(\custom_alu/mult/mult16_3/Q[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[3]_i_5 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[32] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[16] ),
        .O(\custom_alu/mult/mult16_3/Q[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[7]_i_2 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[39] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[23] ),
        .O(\custom_alu/mult/mult16_3/Q[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[7]_i_3 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[38] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[22] ),
        .O(\custom_alu/mult/mult16_3/Q[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[7]_i_4 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[37] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[21] ),
        .O(\custom_alu/mult/mult16_3/Q[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \custom_alu/mult/mult16_3/Q[7]_i_5 
       (.I0(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[36] ),
        .I1(\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[20] ),
        .O(\custom_alu/mult/mult16_3/Q[7]_i_5_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[10]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[27] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[26] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[25] ,\<const0> }),
        .O({\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[10]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[10]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[10]_i_4_n_0 ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[24] }));
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[11]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[43] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[42] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[41] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[40] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[11]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[11]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[11]_i_4_n_0 ,\custom_alu/mult/mult16_3/Q[11]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[14]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[10]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[31] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[30] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[29] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[28] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[14]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[14]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[14]_i_4_n_0 ,\custom_alu/mult/mult16_3/Q[14]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[15]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[11]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[47] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[46] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[45] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[44] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[15]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[15]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[15]_i_4_n_0 ,\custom_alu/mult/mult16_3/Q[15]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[16]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[15]_i_1_n_0 ),
        .CO(\custom_alu/mult/mult16_3/Q_reg[16]_i_1_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const1> }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[18]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[14]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[35] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[34] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[33] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[32] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[18]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[18]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[18]_i_4_n_0 ,\custom_alu/mult/mult16_3/Q[18]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[22]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[18]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[39] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[38] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[37] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[36] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[22]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[22]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[22]_i_4_n_0 ,\custom_alu/mult/mult16_3/Q[22]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[26]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[22]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[41] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[40] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[43] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[42] ,\custom_alu/mult/mult16_3/Q[26]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[26]_i_3_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[30]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[26]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[47] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[46] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[45] ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[44] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[31]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[30]_i_1_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/mult/mult16_3/Q_reg[31]_i_1_n_7 ),
        .S({\<const0> ,\<const0> ,\<const0> ,\custom_alu/mult/mult16_3/FF_MULT_1/Q_reg_n_0_[48] }));
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[35] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[34] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[33] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[32] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[3]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[3]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[3]_i_4_n_0 ,\custom_alu/mult/mult16_3/Q[3]_i_5_n_0 }));
  CARRY4 \custom_alu/mult/mult16_3/Q_reg[7]_i_1 
       (.CI(\custom_alu/mult/mult16_3/Q_reg[3]_i_1_n_0 ),
        .CO({\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_0 ,\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_1 ,\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_2 ,\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[39] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[38] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[37] ,\custom_alu/mult/mult16_3/FF_MULT_0/Q_reg_n_0_[36] }),
        .O({\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_4 ,\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_5 ,\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_6 ,\custom_alu/mult/mult16_3/Q_reg[7]_i_1_n_7 }),
        .S({\custom_alu/mult/mult16_3/Q[7]_i_2_n_0 ,\custom_alu/mult/mult16_3/Q[7]_i_3_n_0 ,\custom_alu/mult/mult16_3/Q[7]_i_4_n_0 ,\custom_alu/mult/mult16_3/Q[7]_i_5_n_0 }));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    exp_b_add_sub_carry__0_i_1
       (.I0(ALU_DIN1[29]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[108]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[29]),
        .O(\custom_alu/fp32_add/p_0_in2_in [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    exp_b_add_sub_carry__0_i_2
       (.I0(ALU_DIN1[28]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[107]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(EX_RF_RD2[28]),
        .O(\custom_alu/fp32_add/p_0_in2_in [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    exp_b_add_sub_carry__0_i_3
       (.I0(ALU_DIN1[27]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[106]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[27]),
        .O(\custom_alu/fp32_add/p_0_in2_in [4]));
  LUT6 #(
    .INIT(64'h555556A6AAAA56A6)) 
    exp_b_add_sub_carry__0_i_4
       (.I0(\custom_alu/fp32_add/p_1_in__0 [7]),
        .I1(EX_RF_RD2[30]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I3(ID_EX_Q[109]),
        .I4(\custom_alu/fp32_add/op_a2 ),
        .I5(ALU_DIN1[30]),
        .O(exp_b_add_sub_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    exp_b_add_sub_carry__0_i_5
       (.I0(EX_RF_RD2[29]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(ID_EX_Q[108]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[29]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [6]),
        .O(exp_b_add_sub_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    exp_b_add_sub_carry__0_i_6
       (.I0(EX_RF_RD2[28]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(ID_EX_Q[107]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[28]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [5]),
        .O(exp_b_add_sub_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    exp_b_add_sub_carry__0_i_7
       (.I0(EX_RF_RD2[27]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(ID_EX_Q[106]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[27]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [4]),
        .O(exp_b_add_sub_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    exp_b_add_sub_carry_i_1
       (.I0(ALU_DIN1[26]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[105]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[26]),
        .O(\custom_alu/fp32_add/p_0_in2_in [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    exp_b_add_sub_carry_i_2
       (.I0(ALU_DIN1[25]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[104]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(EX_RF_RD2[25]),
        .O(\custom_alu/fp32_add/p_0_in2_in [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    exp_b_add_sub_carry_i_3
       (.I0(ALU_DIN1[24]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[103]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[24]),
        .O(\custom_alu/fp32_add/p_0_in2_in [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    exp_b_add_sub_carry_i_4
       (.I0(ALU_DIN1[23]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ID_EX_Q[102]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I4(EX_RF_RD2[23]),
        .O(\custom_alu/fp32_add/p_0_in2_in [0]));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    exp_b_add_sub_carry_i_5
       (.I0(EX_RF_RD2[26]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(ID_EX_Q[105]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[26]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [3]),
        .O(exp_b_add_sub_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    exp_b_add_sub_carry_i_6
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[25]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [2]),
        .O(exp_b_add_sub_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    exp_b_add_sub_carry_i_7
       (.I0(EX_RF_RD2[24]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(ID_EX_Q[103]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[24]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [1]),
        .O(exp_b_add_sub_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    exp_b_add_sub_carry_i_8
       (.I0(EX_RF_RD2[23]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__2_n_0 ),
        .I2(ID_EX_Q[102]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[23]),
        .I5(\custom_alu/fp32_add/p_1_in__0 [0]),
        .O(exp_b_add_sub_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    exp_diff_carry__0_i_1
       (.I0(ID_EX_Q[108]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[29]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[29]),
        .O(exp_diff_carry__0_i_1_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    exp_diff_carry__0_i_2
       (.I0(ID_EX_Q[107]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[28]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[28]),
        .O(exp_diff_carry__0_i_2_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    exp_diff_carry__0_i_3
       (.I0(ID_EX_Q[106]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[27]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[27]),
        .O(exp_diff_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    exp_diff_carry__0_i_4
       (.I0(ID_EX_Q[156]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[30]),
        .I3(ID_EX_Q[109]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[30]),
        .O(exp_diff_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'hE21D)) 
    exp_diff_carry__0_i_5
       (.I0(EX_RF_RD2[29]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[108]),
        .I3(ALU_DIN1[29]),
        .O(exp_diff_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'hE21D)) 
    exp_diff_carry__0_i_6
       (.I0(EX_RF_RD2[28]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[107]),
        .I3(ALU_DIN1[28]),
        .O(exp_diff_carry__0_i_6_n_0));
  LUT4 #(
    .INIT(16'hE21D)) 
    exp_diff_carry__0_i_7
       (.I0(EX_RF_RD2[27]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[106]),
        .I3(ALU_DIN1[27]),
        .O(exp_diff_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    exp_diff_carry_i_1
       (.I0(ID_EX_Q[105]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[26]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[26]),
        .O(exp_diff_carry_i_1_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    exp_diff_carry_i_2
       (.I0(ID_EX_Q[104]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[25]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[25]),
        .O(exp_diff_carry_i_2_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    exp_diff_carry_i_3
       (.I0(ID_EX_Q[103]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[24]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[24]),
        .O(exp_diff_carry_i_3_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    exp_diff_carry_i_4
       (.I0(ID_EX_Q[102]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(EX_RF_RD2[23]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN1[23]),
        .O(exp_diff_carry_i_4_n_0));
  LUT4 #(
    .INIT(16'hE21D)) 
    exp_diff_carry_i_5
       (.I0(EX_RF_RD2[26]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[105]),
        .I3(ALU_DIN1[26]),
        .O(exp_diff_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'hE21D)) 
    exp_diff_carry_i_6
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(ALU_DIN1[25]),
        .O(exp_diff_carry_i_6_n_0));
  LUT4 #(
    .INIT(16'hE21D)) 
    exp_diff_carry_i_7
       (.I0(EX_RF_RD2[24]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[103]),
        .I3(ALU_DIN1[24]),
        .O(exp_diff_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'hE21D)) 
    exp_diff_carry_i_8
       (.I0(EX_RF_RD2[23]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[102]),
        .I3(ALU_DIN1[23]),
        .O(exp_diff_carry_i_8_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    exp_sub_carry__0_i_1
       (.I0(\custom_alu/fp32_add/exp_a [7]),
        .O(exp_sub_carry__0_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    exp_sub_carry__0_i_2
       (.I0(\custom_alu/fp32_add/exp_a [6]),
        .O(exp_sub_carry__0_i_2_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    exp_sub_carry__0_i_3
       (.I0(\custom_alu/fp32_add/exp_a [5]),
        .O(exp_sub_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h5556555555555555)) 
    exp_sub_carry__0_i_4
       (.I0(\custom_alu/fp32_add/exp_a [4]),
        .I1(exp_sub_carry__0_i_5_n_0),
        .I2(\custom_alu/fp32_add/sel0 [21]),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(exp_sub_carry_i_10_n_0),
        .I5(exp_sub_carry__0_i_6_n_0),
        .O(exp_sub_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    exp_sub_carry__0_i_5
       (.I0(exp_sub_carry__0_i_7_n_0),
        .I1(\custom_alu/fp32_add/sel0 [13]),
        .I2(\custom_alu/fp32_add/sel0 [9]),
        .I3(\custom_alu/fp32_add/sel0 [8]),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(exp_sub_carry__0_i_8_n_0),
        .O(exp_sub_carry__0_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT2 #(
    .INIT(4'h1)) 
    exp_sub_carry__0_i_6
       (.I0(\custom_alu/fp32_add/sel0 [11]),
        .I1(\custom_alu/fp32_add/sel0 [10]),
        .O(exp_sub_carry__0_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    exp_sub_carry__0_i_7
       (.I0(\custom_alu/fp32_add/sel0 [16]),
        .I1(\custom_alu/fp32_add/sel0 [14]),
        .I2(\custom_alu/fp32_add/sel0 [12]),
        .O(exp_sub_carry__0_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    exp_sub_carry__0_i_8
       (.I0(\custom_alu/fp32_add/sel0 [18]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [20]),
        .I3(\custom_alu/fp32_add/sel0 [19]),
        .O(exp_sub_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h6555666666666666)) 
    exp_sub_carry_i_1
       (.I0(\custom_alu/fp32_add/exp_a [3]),
        .I1(exp_sub_carry_i_5_n_0),
        .I2(exp_sub_carry_i_6_n_0),
        .I3(exp_sub_carry_i_7_n_0),
        .I4(exp_sub_carry_i_8_n_0),
        .I5(exp_sub_carry_i_9_n_0),
        .O(exp_sub_carry_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT2 #(
    .INIT(4'h2)) 
    exp_sub_carry_i_10
       (.I0(\custom_alu/fp32_add/sel0 [24]),
        .I1(\custom_alu/fp32_add/sel0 [23]),
        .O(exp_sub_carry_i_10_n_0));
  LUT6 #(
    .INIT(64'h0001000000010001)) 
    exp_sub_carry_i_11
       (.I0(\custom_alu/fp32_add/sel0 [16]),
        .I1(\custom_alu/fp32_add/sel0 [17]),
        .I2(\custom_alu/fp32_add/sel0 [18]),
        .I3(\custom_alu/fp32_add/sel0 [19]),
        .I4(exp_sub_carry_i_17_n_0),
        .I5(exp_sub_carry_i_8_n_0),
        .O(exp_sub_carry_i_11_n_0));
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT2 #(
    .INIT(4'h1)) 
    exp_sub_carry_i_12
       (.I0(\custom_alu/fp32_add/sel0 [21]),
        .I1(\custom_alu/fp32_add/sel0 [20]),
        .O(exp_sub_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h1111111111110010)) 
    exp_sub_carry_i_13
       (.I0(\custom_alu/fp32_add/sel0 [17]),
        .I1(\custom_alu/fp32_add/sel0 [16]),
        .I2(exp_sub_carry_i_18_n_0),
        .I3(exp_sub_carry_i_19_n_0),
        .I4(\custom_alu/fp32_add/sel0 [15]),
        .I5(\custom_alu/fp32_add/sel0 [14]),
        .O(exp_sub_carry_i_13_n_0));
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT2 #(
    .INIT(4'h1)) 
    exp_sub_carry_i_14
       (.I0(\custom_alu/fp32_add/sel0 [18]),
        .I1(\custom_alu/fp32_add/sel0 [19]),
        .O(exp_sub_carry_i_14_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00AB)) 
    exp_sub_carry_i_15
       (.I0(\custom_alu/fp32_add/sel0 [19]),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(exp_sub_carry_i_20_n_0),
        .I3(\custom_alu/fp32_add/sel0 [20]),
        .I4(\custom_alu/fp32_add/sel0 [21]),
        .I5(\custom_alu/fp32_add/sel0 [22]),
        .O(exp_sub_carry_i_15_n_0));
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT4 #(
    .INIT(16'hFFFB)) 
    exp_sub_carry_i_16
       (.I0(\custom_alu/fp32_add/sel0 [23]),
        .I1(\custom_alu/fp32_add/sel0 [24]),
        .I2(\custom_alu/fp32_add/sel0 [22]),
        .I3(\custom_alu/fp32_add/sel0 [21]),
        .O(exp_sub_carry_i_16_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    exp_sub_carry_i_17
       (.I0(exp_sub_carry_i_9_n_0),
        .I1(exp_sub_carry_i_6_n_0),
        .I2(\custom_alu/fp32_add/sel0 [4]),
        .I3(\custom_alu/fp32_add/sel0 [5]),
        .I4(\custom_alu/fp32_add/sel0 [7]),
        .I5(\custom_alu/fp32_add/sel0 [6]),
        .O(exp_sub_carry_i_17_n_0));
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT2 #(
    .INIT(4'h1)) 
    exp_sub_carry_i_18
       (.I0(\custom_alu/fp32_add/sel0 [12]),
        .I1(\custom_alu/fp32_add/sel0 [13]),
        .O(exp_sub_carry_i_18_n_0));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8A8A8AA)) 
    exp_sub_carry_i_19
       (.I0(exp_sub_carry__0_i_6_n_0),
        .I1(\custom_alu/fp32_add/sel0 [8]),
        .I2(\custom_alu/fp32_add/sel0 [9]),
        .I3(\custom_alu/fp32_add/sel0 [7]),
        .I4(\custom_alu/fp32_add/sel0 [6]),
        .I5(exp_sub_carry_i_21_n_0),
        .O(exp_sub_carry_i_19_n_0));
  LUT6 #(
    .INIT(64'h5555555555565555)) 
    exp_sub_carry_i_2
       (.I0(\custom_alu/fp32_add/exp_a [2]),
        .I1(\custom_alu/fp32_add/sel0 [20]),
        .I2(\custom_alu/fp32_add/sel0 [21]),
        .I3(\custom_alu/fp32_add/sel0 [22]),
        .I4(exp_sub_carry_i_10_n_0),
        .I5(exp_sub_carry_i_11_n_0),
        .O(exp_sub_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h88A888AA88A888A8)) 
    exp_sub_carry_i_20
       (.I0(exp_sub_carry_i_22_n_0),
        .I1(exp_sub_carry__0_i_7_n_0),
        .I2(\custom_alu/fp32_add/sel0 [10]),
        .I3(\custom_alu/fp32_add/sel0 [11]),
        .I4(\custom_alu/fp32_add/sel0 [9]),
        .I5(exp_sub_carry_i_23_n_0),
        .O(exp_sub_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'h1110111011101111)) 
    exp_sub_carry_i_21
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [5]),
        .I2(\custom_alu/fp32_add/sel0 [2]),
        .I3(\custom_alu/fp32_add/sel0 [3]),
        .I4(\custom_alu/fp32_add/sel0 [1]),
        .I5(\custom_alu/fp32_add/sel0 [0]),
        .O(exp_sub_carry_i_21_n_0));
  LUT5 #(
    .INIT(32'h0000FF0D)) 
    exp_sub_carry_i_22
       (.I0(\custom_alu/fp32_add/sel0 [13]),
        .I1(\custom_alu/fp32_add/sel0 [14]),
        .I2(\custom_alu/fp32_add/sel0 [15]),
        .I3(\custom_alu/fp32_add/sel0 [16]),
        .I4(\custom_alu/fp32_add/sel0 [17]),
        .O(exp_sub_carry_i_22_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFEFEE)) 
    exp_sub_carry_i_23
       (.I0(\custom_alu/fp32_add/sel0 [8]),
        .I1(\custom_alu/fp32_add/sel0 [6]),
        .I2(\custom_alu/fp32_add/sel0 [5]),
        .I3(\custom_alu/fp32_add/sel0 [4]),
        .I4(exp_sub_carry_i_24_n_0),
        .I5(\custom_alu/fp32_add/sel0 [7]),
        .O(exp_sub_carry_i_23_n_0));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT5 #(
    .INIT(32'h000000F2)) 
    exp_sub_carry_i_24
       (.I0(\custom_alu/fp32_add/sel0 [0]),
        .I1(\custom_alu/fp32_add/sel0 [1]),
        .I2(\custom_alu/fp32_add/sel0 [2]),
        .I3(\custom_alu/fp32_add/sel0 [3]),
        .I4(\custom_alu/fp32_add/sel0 [5]),
        .O(exp_sub_carry_i_24_n_0));
  LUT6 #(
    .INIT(64'h5565656555655565)) 
    exp_sub_carry_i_3
       (.I0(\custom_alu/fp32_add/exp_a [1]),
        .I1(\custom_alu/fp32_add/sel0 [22]),
        .I2(exp_sub_carry_i_10_n_0),
        .I3(exp_sub_carry_i_12_n_0),
        .I4(exp_sub_carry_i_13_n_0),
        .I5(exp_sub_carry_i_14_n_0),
        .O(exp_sub_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h5559)) 
    exp_sub_carry_i_4
       (.I0(\custom_alu/fp32_add/exp_a [0]),
        .I1(\custom_alu/fp32_add/sel0 [24]),
        .I2(\custom_alu/fp32_add/sel0 [23]),
        .I3(exp_sub_carry_i_15_n_0),
        .O(exp_sub_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    exp_sub_carry_i_5
       (.I0(exp_sub_carry_i_16_n_0),
        .I1(\custom_alu/fp32_add/sel0 [18]),
        .I2(\custom_alu/fp32_add/sel0 [17]),
        .I3(\custom_alu/fp32_add/sel0 [20]),
        .I4(\custom_alu/fp32_add/sel0 [19]),
        .I5(\custom_alu/fp32_add/sel0 [16]),
        .O(exp_sub_carry_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    exp_sub_carry_i_6
       (.I0(\custom_alu/fp32_add/sel0 [0]),
        .I1(\custom_alu/fp32_add/sel0 [1]),
        .I2(\custom_alu/fp32_add/sel0 [3]),
        .I3(\custom_alu/fp32_add/sel0 [2]),
        .O(exp_sub_carry_i_6_n_0));
  LUT4 #(
    .INIT(16'h0001)) 
    exp_sub_carry_i_7
       (.I0(\custom_alu/fp32_add/sel0 [4]),
        .I1(\custom_alu/fp32_add/sel0 [5]),
        .I2(\custom_alu/fp32_add/sel0 [7]),
        .I3(\custom_alu/fp32_add/sel0 [6]),
        .O(exp_sub_carry_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    exp_sub_carry_i_8
       (.I0(\custom_alu/fp32_add/sel0 [13]),
        .I1(\custom_alu/fp32_add/sel0 [12]),
        .I2(\custom_alu/fp32_add/sel0 [14]),
        .I3(\custom_alu/fp32_add/sel0 [15]),
        .O(exp_sub_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h0001)) 
    exp_sub_carry_i_9
       (.I0(\custom_alu/fp32_add/sel0 [10]),
        .I1(\custom_alu/fp32_add/sel0 [11]),
        .I2(\custom_alu/fp32_add/sel0 [9]),
        .I3(\custom_alu/fp32_add/sel0 [8]),
        .O(exp_sub_carry_i_9_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    exponent_carry__0_i_1
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[62] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[30] ),
        .O(exponent_carry__0_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    exponent_carry__0_i_2
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[28] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[60] ),
        .O(exponent_carry__0_i_2_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    exponent_carry__0_i_3
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[27] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[59] ),
        .O(exponent_carry__0_i_3_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    exponent_carry__0_i_4
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[26] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[58] ),
        .O(exponent_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h6999)) 
    exponent_carry__0_i_5
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[30] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[62] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[61] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[29] ),
        .O(exponent_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    exponent_carry__0_i_6
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[60] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[28] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[61] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[29] ),
        .O(exponent_carry__0_i_6_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    exponent_carry__0_i_7
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[59] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[27] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[60] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[28] ),
        .O(exponent_carry__0_i_7_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    exponent_carry__0_i_8
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[58] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[26] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[59] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[27] ),
        .O(exponent_carry__0_i_8_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    exponent_carry__1_i_1
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[30] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[62] ),
        .O(exponent_carry__1_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    exponent_carry_i_1
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[25] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[57] ),
        .O(exponent_carry_i_1_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 exponent_carry_i_10
       (.CI(exponent_carry_i_11_n_0),
        .CO({exponent_carry_i_10_n_0,exponent_carry_i_10_n_1,exponent_carry_i_10_n_2,exponent_carry_i_10_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({exponent_carry_i_10_n_4,exponent_carry_i_10_n_5,exponent_carry_i_10_n_6,exponent_carry_i_10_n_7}),
        .S(\custom_alu/fp32_mult/p_1_in [42:39]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 exponent_carry_i_11
       (.CI(\Q_reg[16]_i_13_n_0 ),
        .CO({exponent_carry_i_11_n_0,exponent_carry_i_11_n_1,exponent_carry_i_11_n_2,exponent_carry_i_11_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\custom_alu/fp32_mult/p_1_in [36:35]}),
        .O({exponent_carry_i_11_n_4,exponent_carry_i_11_n_5,exponent_carry_i_11_n_6,exponent_carry_i_11_n_7}),
        .S({\custom_alu/fp32_mult/p_1_in [38:37],\fp32_mult/mult24_0/exponent_carry_i_12_n_0 ,\fp32_mult/mult24_0/exponent_carry_i_13_n_0 }));
  LUT2 #(
    .INIT(4'h8)) 
    exponent_carry_i_2
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[24] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[56] ),
        .O(exponent_carry_i_2_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    exponent_carry_i_3
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[23] ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .O(exponent_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    exponent_carry_i_4
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[57] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[25] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[58] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[26] ),
        .O(exponent_carry_i_4_n_0));
  LUT4 #(
    .INIT(16'h8778)) 
    exponent_carry_i_5
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[56] ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[24] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[57] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[25] ),
        .O(exponent_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'hE11E)) 
    exponent_carry_i_6
       (.I0(\custom_alu/fp32_mult/normalised ),
        .I1(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[23] ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[56] ),
        .I3(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[24] ),
        .O(exponent_carry_i_6_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    exponent_carry_i_7
       (.I0(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[23] ),
        .I1(\custom_alu/fp32_mult/normalised ),
        .I2(\custom_alu/fp32_mult/FF_MULT_2/Q_reg_n_0_[55] ),
        .O(exponent_carry_i_7_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 exponent_carry_i_8
       (.CI(exponent_carry_i_9_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\custom_alu/fp32_mult/normalised ),
        .S({\<const0> ,\<const0> ,\<const0> ,\custom_alu/fp32_mult/p_1_in [47]}));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 exponent_carry_i_9
       (.CI(exponent_carry_i_10_n_0),
        .CO({exponent_carry_i_9_n_0,exponent_carry_i_9_n_1,exponent_carry_i_9_n_2,exponent_carry_i_9_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({exponent_carry_i_9_n_4,exponent_carry_i_9_n_5,exponent_carry_i_9_n_6,exponent_carry_i_9_n_7}),
        .S(\custom_alu/fp32_mult/p_1_in [46:43]));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[12]_i_10 
       (.I0(ALU_DIN1[8]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[8]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[87]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [8]),
        .O(\fp32_add/Q[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[12]_i_7 
       (.I0(ALU_DIN1[11]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[11]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[90]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [11]),
        .O(\fp32_add/Q[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[12]_i_8 
       (.I0(ALU_DIN1[10]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[10]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[89]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [10]),
        .O(\fp32_add/Q[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[12]_i_9 
       (.I0(ALU_DIN1[9]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[9]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[88]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [9]),
        .O(\fp32_add/Q[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[16]_i_10 
       (.I0(ALU_DIN1[12]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[12]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[91]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [12]),
        .O(\fp32_add/Q[16]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[16]_i_7 
       (.I0(ALU_DIN1[15]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[15]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[94]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [15]),
        .O(\fp32_add/Q[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[16]_i_8 
       (.I0(ALU_DIN1[14]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[14]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[93]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [14]),
        .O(\fp32_add/Q[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[16]_i_9 
       (.I0(ALU_DIN1[13]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[13]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[92]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [13]),
        .O(\fp32_add/Q[16]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h9A999AAA)) 
    \fp32_add/Q[20]_i_10 
       (.I0(\Q[20]_i_18_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[20]_i_13__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_14__1_n_0 ),
        .O(\fp32_add/Q[20]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h9A999AAA)) 
    \fp32_add/Q[20]_i_7 
       (.I0(\Q[20]_i_15_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[23]_i_15_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_11__1_n_0 ),
        .O(\fp32_add/Q[20]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h9A999AAA)) 
    \fp32_add/Q[20]_i_8 
       (.I0(\Q[20]_i_16_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[20]_i_11__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_12__1_n_0 ),
        .O(\fp32_add/Q[20]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h9A999AAA)) 
    \fp32_add/Q[20]_i_9 
       (.I0(\Q[20]_i_17_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[20]_i_12__1_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[20]_i_13__1_n_0 ),
        .O(\fp32_add/Q[20]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h9A999AAA)) 
    \fp32_add/Q[23]_i_10 
       (.I0(\Q[23]_i_17_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[23]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[23]_i_15_n_0 ),
        .O(\fp32_add/Q[23]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[23]_i_8 
       (.I0(ALU_DIN1[22]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[22]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[101]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [22]),
        .O(\fp32_add/Q[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAA9A9999AA9AAAAA)) 
    \fp32_add/Q[23]_i_9 
       (.I0(\Q[23]_i_16_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[23]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [1]),
        .I4(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I5(\Q[23]_i_14_n_0 ),
        .O(\fp32_add/Q[23]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E21DE21DE21D)) 
    \fp32_add/Q[4]_i_10 
       (.I0(ALU_DIN1[0]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(ALU_DIN2[0]),
        .I3(\Q[4]_i_19_n_0 ),
        .I4(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I5(\Q[4]_i_13_n_0 ),
        .O(\fp32_add/Q[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h9AAA9A99)) 
    \fp32_add/Q[4]_i_7 
       (.I0(\Q[4]_i_16_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[8]_i_14_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[4]_i_11_n_0 ),
        .O(\fp32_add/Q[4]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hAA9A999A)) 
    \fp32_add/Q[4]_i_8 
       (.I0(\Q[4]_i_17_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[4]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[4]_i_11_n_0 ),
        .O(\fp32_add/Q[4]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h9AAA9A99)) 
    \fp32_add/Q[4]_i_9 
       (.I0(\Q[4]_i_18_n_0 ),
        .I1(\Q[23]_i_13_n_0 ),
        .I2(\Q[4]_i_12_n_0 ),
        .I3(\custom_alu/fp32_add/p_1_in__0 [0]),
        .I4(\Q[4]_i_13_n_0 ),
        .O(\fp32_add/Q[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[67]_i_4 
       (.I0(EX_RF_RD1[3]),
        .I1(\FF_ID_EX/Q_reg_n_0_[170] ),
        .I2(ID_EX_Q[129]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN2[3]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [3]),
        .O(\fp32_add/Q[67]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[67]_i_5 
       (.I0(EX_RF_RD1[2]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[128]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN2[2]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [2]),
        .O(\fp32_add/Q[67]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[67]_i_6 
       (.I0(EX_RF_RD1[1]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[127]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN2[1]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [1]),
        .O(\fp32_add/Q[67]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[67]_i_7 
       (.I0(EX_RF_RD1[0]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[126]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN2[0]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [0]),
        .O(\fp32_add/Q[67]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[71]_i_4 
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[7]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[86]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [7]),
        .O(\fp32_add/Q[71]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[71]_i_5 
       (.I0(ALU_DIN1[6]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[6]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[85]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [6]),
        .O(\fp32_add/Q[71]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[71]_i_6 
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN2[5]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [5]),
        .O(\fp32_add/Q[71]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[71]_i_7 
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(op_a2_carry_i_9_n_0),
        .I5(\custom_alu/fp32_add/significand_sub_complement [4]),
        .O(\fp32_add/Q[71]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[75]_i_4 
       (.I0(ALU_DIN1[11]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[11]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[90]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [11]),
        .O(\fp32_add/Q[75]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[75]_i_5 
       (.I0(ALU_DIN1[10]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[10]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[89]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [10]),
        .O(\fp32_add/Q[75]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[75]_i_6 
       (.I0(ALU_DIN1[9]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[9]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[88]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [9]),
        .O(\fp32_add/Q[75]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[75]_i_7 
       (.I0(ALU_DIN1[8]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[8]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[87]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [8]),
        .O(\fp32_add/Q[75]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[79]_i_4 
       (.I0(ALU_DIN1[15]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[15]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[94]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [15]),
        .O(\fp32_add/Q[79]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[79]_i_5 
       (.I0(ALU_DIN1[14]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[14]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[93]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [14]),
        .O(\fp32_add/Q[79]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[79]_i_6 
       (.I0(ALU_DIN1[13]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[13]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[92]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [13]),
        .O(\fp32_add/Q[79]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[79]_i_7 
       (.I0(ALU_DIN1[12]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[12]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[91]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [12]),
        .O(\fp32_add/Q[79]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[83]_i_4 
       (.I0(ALU_DIN1[19]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[19]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[98]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [19]),
        .O(\fp32_add/Q[83]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[83]_i_5 
       (.I0(ALU_DIN1[18]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[18]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[97]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [18]),
        .O(\fp32_add/Q[83]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[83]_i_6 
       (.I0(ALU_DIN1[17]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[17]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[96]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [17]),
        .O(\fp32_add/Q[83]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[83]_i_7 
       (.I0(ALU_DIN1[16]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[16]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[95]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [16]),
        .O(\fp32_add/Q[83]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[87]_i_5 
       (.I0(ALU_DIN1[22]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[22]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[101]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [22]),
        .O(\fp32_add/Q[87]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[87]_i_6 
       (.I0(ALU_DIN1[21]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[21]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[100]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [21]),
        .O(\fp32_add/Q[87]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[87]_i_7 
       (.I0(ALU_DIN1[20]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[20]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[99]),
        .I5(\custom_alu/fp32_add/significand_sub_complement [20]),
        .O(\fp32_add/Q[87]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[8]_i_10 
       (.I0(EX_RF_RD1[4]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[130]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(op_a2_carry_i_9_n_0),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [4]),
        .O(\fp32_add/Q[8]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[8]_i_7 
       (.I0(ALU_DIN1[7]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[7]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[86]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [7]),
        .O(\fp32_add/Q[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DEEE222E2)) 
    \fp32_add/Q[8]_i_8 
       (.I0(ALU_DIN1[6]),
        .I1(\custom_alu/fp32_add/op_a2 ),
        .I2(EX_RF_RD2[6]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I4(ID_EX_Q[85]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [6]),
        .O(\fp32_add/Q[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \fp32_add/Q[8]_i_9 
       (.I0(EX_RF_RD1[5]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(ID_EX_Q[131]),
        .I3(\custom_alu/fp32_add/op_a2 ),
        .I4(ALU_DIN2[5]),
        .I5(\custom_alu/fp32_add/significand_b_add_sub [5]),
        .O(\fp32_add/Q[8]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[16]_i_14 
       (.I0(\custom_alu/fp32_mult/p_1_in [34]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[22] ),
        .O(\fp32_mult/mult24_0/Q[16]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[16]_i_15 
       (.I0(\custom_alu/fp32_mult/p_1_in [33]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[21] ),
        .O(\fp32_mult/mult24_0/Q[16]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[16]_i_16 
       (.I0(\custom_alu/fp32_mult/p_1_in [32]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[20] ),
        .O(\fp32_mult/mult24_0/Q[16]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[16]_i_17 
       (.I0(\custom_alu/fp32_mult/p_1_in [31]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[19] ),
        .O(\fp32_mult/mult24_0/Q[16]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_24 
       (.I0(\custom_alu/fp32_mult/p_1_in [26]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[14] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_25 
       (.I0(\custom_alu/fp32_mult/p_1_in [25]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[13] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_26 
       (.I0(\custom_alu/fp32_mult/p_1_in [24]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[12] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_27 
       (.I0(\custom_alu/fp32_mult/p_1_in [23]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[11] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_28 
       (.I0(\custom_alu/fp32_mult/p_1_in [30]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[18] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_29 
       (.I0(\custom_alu/fp32_mult/p_1_in [29]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[17] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_30 
       (.I0(\custom_alu/fp32_mult/p_1_in [28]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[16] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_31 
       (.I0(\custom_alu/fp32_mult/p_1_in [27]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[15] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_37 
       (.I0(\custom_alu/fp32_mult/p_1_in [22]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[10] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_37_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_38 
       (.I0(\custom_alu/fp32_mult/p_1_in [21]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[9] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_39 
       (.I0(\custom_alu/fp32_mult/p_1_in [20]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[8] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_39_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_40 
       (.I0(\custom_alu/fp32_mult/p_1_in [19]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[7] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_41 
       (.I0(\custom_alu/fp32_mult/p_1_in [14]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[2] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_42 
       (.I0(\custom_alu/fp32_mult/p_1_in [13]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[1] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_43 
       (.I0(\custom_alu/fp32_mult/p_1_in [12]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[0] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_43_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_44 
       (.I0(\custom_alu/fp32_mult/p_1_in [18]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[6] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_45 
       (.I0(\custom_alu/fp32_mult/p_1_in [17]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[5] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_46 
       (.I0(\custom_alu/fp32_mult/p_1_in [16]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[4] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/Q[49]_i_47 
       (.I0(\custom_alu/fp32_mult/p_1_in [15]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[3] ),
        .O(\fp32_mult/mult24_0/Q[49]_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/exponent_carry_i_12 
       (.I0(\custom_alu/fp32_mult/p_1_in [36]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[24] ),
        .O(\fp32_mult/mult24_0/exponent_carry_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \fp32_mult/mult24_0/exponent_carry_i_13 
       (.I0(\custom_alu/fp32_mult/p_1_in [35]),
        .I1(\custom_alu/fp32_mult/mult24_0/FF_MULT_1/Q_reg_n_0_[23] ),
        .O(\fp32_mult/mult24_0/exponent_carry_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__0_i_1
       (.I0(ALU_DIN2[15]),
        .I1(ALU_DIN1[15]),
        .I2(EX_RF_RD2[14]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[93]),
        .I5(ALU_DIN1[14]),
        .O(op_a2_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__0_i_2
       (.I0(ALU_DIN2[13]),
        .I1(ALU_DIN1[13]),
        .I2(EX_RF_RD2[12]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[91]),
        .I5(ALU_DIN1[12]),
        .O(op_a2_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__0_i_3
       (.I0(ALU_DIN2[11]),
        .I1(ALU_DIN1[11]),
        .I2(EX_RF_RD2[10]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[89]),
        .I5(ALU_DIN1[10]),
        .O(op_a2_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'h00E200E2E2FF00E2)) 
    op_a2_carry__0_i_4
       (.I0(EX_RF_RD2[9]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[88]),
        .I3(ALU_DIN1[9]),
        .I4(ALU_DIN2[8]),
        .I5(ALU_DIN1[8]),
        .O(op_a2_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__0_i_5
       (.I0(ALU_DIN1[15]),
        .I1(ID_EX_Q[94]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[15]),
        .I4(ALU_DIN1[14]),
        .I5(ALU_DIN2[14]),
        .O(op_a2_carry__0_i_5_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__0_i_6
       (.I0(ALU_DIN1[13]),
        .I1(ID_EX_Q[92]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[13]),
        .I4(ALU_DIN1[12]),
        .I5(ALU_DIN2[12]),
        .O(op_a2_carry__0_i_6_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__0_i_7
       (.I0(ALU_DIN1[11]),
        .I1(ID_EX_Q[90]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[11]),
        .I4(ALU_DIN1[10]),
        .I5(ALU_DIN2[10]),
        .O(op_a2_carry__0_i_7_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__0_i_8
       (.I0(ALU_DIN1[9]),
        .I1(ID_EX_Q[88]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[9]),
        .I4(ALU_DIN1[8]),
        .I5(ALU_DIN2[8]),
        .O(op_a2_carry__0_i_8_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__1_i_1
       (.I0(ALU_DIN2[23]),
        .I1(ALU_DIN1[23]),
        .I2(EX_RF_RD2[22]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[101]),
        .I5(ALU_DIN1[22]),
        .O(op_a2_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__1_i_2
       (.I0(ALU_DIN2[21]),
        .I1(ALU_DIN1[21]),
        .I2(EX_RF_RD2[20]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[99]),
        .I5(ALU_DIN1[20]),
        .O(op_a2_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__1_i_3
       (.I0(ALU_DIN2[19]),
        .I1(ALU_DIN1[19]),
        .I2(EX_RF_RD2[18]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[97]),
        .I5(ALU_DIN1[18]),
        .O(op_a2_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'h00E200E2E2FF00E2)) 
    op_a2_carry__1_i_4
       (.I0(EX_RF_RD2[17]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[96]),
        .I3(ALU_DIN1[17]),
        .I4(ALU_DIN2[16]),
        .I5(ALU_DIN1[16]),
        .O(op_a2_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__1_i_5
       (.I0(ALU_DIN1[23]),
        .I1(ID_EX_Q[102]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(EX_RF_RD2[23]),
        .I4(ALU_DIN1[22]),
        .I5(ALU_DIN2[22]),
        .O(op_a2_carry__1_i_5_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__1_i_6
       (.I0(ALU_DIN1[21]),
        .I1(ID_EX_Q[100]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(EX_RF_RD2[21]),
        .I4(ALU_DIN1[20]),
        .I5(ALU_DIN2[20]),
        .O(op_a2_carry__1_i_6_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__1_i_7
       (.I0(ALU_DIN1[19]),
        .I1(ID_EX_Q[98]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(EX_RF_RD2[19]),
        .I4(ALU_DIN1[18]),
        .I5(ALU_DIN2[18]),
        .O(op_a2_carry__1_i_7_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__1_i_8
       (.I0(ALU_DIN1[17]),
        .I1(ID_EX_Q[96]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[17]),
        .I4(ALU_DIN1[16]),
        .I5(ALU_DIN2[16]),
        .O(op_a2_carry__1_i_8_n_0));
  LUT6 #(
    .INIT(64'h000000E2E2E200E2)) 
    op_a2_carry__2_i_1
       (.I0(EX_RF_RD2[30]),
        .I1(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I2(ID_EX_Q[109]),
        .I3(EX_RF_RD1[30]),
        .I4(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I5(ID_EX_Q[156]),
        .O(op_a2_carry__2_i_1_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__2_i_2
       (.I0(ALU_DIN2[29]),
        .I1(ALU_DIN1[29]),
        .I2(EX_RF_RD2[28]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[107]),
        .I5(ALU_DIN1[28]),
        .O(op_a2_carry__2_i_2_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry__2_i_3
       (.I0(ALU_DIN2[27]),
        .I1(ALU_DIN1[27]),
        .I2(EX_RF_RD2[26]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[105]),
        .I5(ALU_DIN1[26]),
        .O(op_a2_carry__2_i_3_n_0));
  LUT6 #(
    .INIT(64'h00E200E2E2FF00E2)) 
    op_a2_carry__2_i_4
       (.I0(EX_RF_RD2[25]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(ID_EX_Q[104]),
        .I3(ALU_DIN1[25]),
        .I4(ALU_DIN2[24]),
        .I5(ALU_DIN1[24]),
        .O(op_a2_carry__2_i_4_n_0));
  LUT6 #(
    .INIT(64'hB847B8B8B8474747)) 
    op_a2_carry__2_i_5
       (.I0(ID_EX_Q[156]),
        .I1(\FF_ID_EX/Q_reg[170]_rep_n_0 ),
        .I2(EX_RF_RD1[30]),
        .I3(ID_EX_Q[109]),
        .I4(\FF_ID_EX/Q_reg[158]_rep_n_0 ),
        .I5(EX_RF_RD2[30]),
        .O(op_a2_carry__2_i_5_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__2_i_6
       (.I0(ALU_DIN1[29]),
        .I1(ID_EX_Q[108]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(EX_RF_RD2[29]),
        .I4(ALU_DIN1[28]),
        .I5(ALU_DIN2[28]),
        .O(op_a2_carry__2_i_6_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__2_i_7
       (.I0(ALU_DIN1[27]),
        .I1(ID_EX_Q[106]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__4_n_0 ),
        .I3(EX_RF_RD2[27]),
        .I4(ALU_DIN1[26]),
        .I5(ALU_DIN2[26]),
        .O(op_a2_carry__2_i_7_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry__2_i_8
       (.I0(ALU_DIN1[25]),
        .I1(ID_EX_Q[104]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[25]),
        .I4(ALU_DIN1[24]),
        .I5(ALU_DIN2[24]),
        .O(op_a2_carry__2_i_8_n_0));
  LUT6 #(
    .INIT(64'h22222222BBB222B2)) 
    op_a2_carry_i_1
       (.I0(ALU_DIN2[7]),
        .I1(ALU_DIN1[7]),
        .I2(EX_RF_RD2[6]),
        .I3(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I4(ID_EX_Q[85]),
        .I5(ALU_DIN1[6]),
        .O(op_a2_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    op_a2_carry_i_2
       (.I0(ALU_DIN2[5]),
        .I1(ALU_DIN1[5]),
        .I2(op_a2_carry_i_9_n_0),
        .I3(EX_RF_RD1[4]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I5(ID_EX_Q[130]),
        .O(op_a2_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    op_a2_carry_i_3
       (.I0(ALU_DIN2[3]),
        .I1(ALU_DIN1[3]),
        .I2(ALU_DIN2[2]),
        .I3(EX_RF_RD1[2]),
        .I4(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I5(ID_EX_Q[128]),
        .O(op_a2_carry_i_3_n_0));
  LUT6 #(
    .INIT(64'h02A202A2ABFB02A2)) 
    op_a2_carry_i_4
       (.I0(ALU_DIN2[1]),
        .I1(EX_RF_RD1[1]),
        .I2(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I3(ID_EX_Q[127]),
        .I4(ALU_DIN2[0]),
        .I5(ALU_DIN1[0]),
        .O(op_a2_carry_i_4_n_0));
  LUT6 #(
    .INIT(64'h9A95000000009A95)) 
    op_a2_carry_i_5
       (.I0(ALU_DIN1[7]),
        .I1(ID_EX_Q[86]),
        .I2(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I3(EX_RF_RD2[7]),
        .I4(ALU_DIN1[6]),
        .I5(ALU_DIN2[6]),
        .O(op_a2_carry_i_5_n_0));
  LUT6 #(
    .INIT(64'h9099900009000999)) 
    op_a2_carry_i_6
       (.I0(ALU_DIN1[5]),
        .I1(ALU_DIN2[5]),
        .I2(ID_EX_Q[130]),
        .I3(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I4(EX_RF_RD1[4]),
        .I5(op_a2_carry_i_9_n_0),
        .O(op_a2_carry_i_6_n_0));
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    op_a2_carry_i_7
       (.I0(ID_EX_Q[129]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[3]),
        .I3(ALU_DIN2[3]),
        .I4(ALU_DIN1[2]),
        .I5(ALU_DIN2[2]),
        .O(op_a2_carry_i_7_n_0));
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    op_a2_carry_i_8
       (.I0(ID_EX_Q[127]),
        .I1(\FF_ID_EX/Q_reg[170]_rep__3_n_0 ),
        .I2(EX_RF_RD1[1]),
        .I3(ALU_DIN2[1]),
        .I4(ALU_DIN1[0]),
        .I5(ALU_DIN2[0]),
        .O(op_a2_carry_i_8_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    op_a2_carry_i_9
       (.I0(ID_EX_Q[83]),
        .I1(\FF_ID_EX/Q_reg[158]_rep__3_n_0 ),
        .I2(EX_RF_RD2[4]),
        .O(op_a2_carry_i_9_n_0));
endmodule
